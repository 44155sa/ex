module TEMAC_CORE_df9b4c715b25(reset, mac_has_sgmii, rx_correct_frame, rx_error_frame, rx_data, rx_data_vld, rx_status_vector, rx_status_vld, rx_clk_en, tx_data, tx_data_en, tx_stop, tx_rdy, tx_retransmit, tx_collision, tx_clk_en, tx_ifg_val, tx_status_vector, tx_status_vld, pause_req, pause_val,
tx_mac_clk, rx_mac_clk, speed_1000,speed_100, speed_10, gmii_col, gmii_crs, gmii_tx_clken, gmii_txd, gmii_tx_en, gmii_tx_er, gmii_rxd, gmii_rx_vld, gmii_rx_er, mdio_in, mdio_out, mdio_oen, mdio_clk,
s_axi_aclk, s_axi_awaddr, s_axi_awvalid, s_axi_awready, s_axi_wdata, s_axi_wvalid, s_axi_wready, s_axi_bresp, s_axi_bvalid, s_axi_bready, s_axi_araddr, s_axi_arvalid, s_axi_arready, s_axi_rdata, s_axi_rresp, s_axi_rvalid, s_axi_rready,
mac_cfg_vector, unicast_addr,pause_source_addr,
ptp_timer_format_i, tx_1588v2_cmd_i, tx_system_time_i, tx_timestamp_i, tx_timestamp_o, tx_tagid_o, tx_timestamp_valid_o, tx_1588v2_cfg_err_o, rx_phy_timer_i, rx_timestamp_o, rx_timestamp_valid_o);
parameter     P_HALF_DUPLEX 	    = 1'b0;		
parameter     P_HOST_EN 	        = 1'b0;		
parameter     P_ADD_FILT_EN 	    = 1'b1;     
parameter     P_ADD_FILT_LIST 	= 0;		
parameter     P_SPEED_10_100     = 1'b0;		
parameter     P_SPEED_1000 	    = 1'b0;		
parameter     P_TRI_SPEED 	    = 1'b1;		
parameter     CFG_1588V2         = 1'b0;   	
input         reset;
input         tx_mac_clk;
input         rx_mac_clk;
output        speed_1000;
output        speed_100;
output        speed_10;
input		 mac_has_sgmii;
input         tx_clk_en;
input  [7:0]  tx_data;
input         tx_data_en;
output        tx_rdy;
input         tx_stop;
output        tx_retransmit;
output        tx_collision;
input  [7:0]  tx_ifg_val;
output [28:0] tx_status_vector;
output        tx_status_vld;
input         rx_clk_en;
output [7:0]  rx_data;
output        rx_data_vld;
output        rx_correct_frame;
output        rx_error_frame;
output [26:0] rx_status_vector;
output        rx_status_vld;
input         pause_req;
input [15:0]  pause_val;
input [47:0]  pause_source_addr;
input [47:0]  unicast_addr;
input          s_axi_aclk;
input  [7 : 0] s_axi_awaddr;
input          s_axi_awvalid;
output         s_axi_awready;
input  [31: 0] s_axi_wdata;
input          s_axi_wvalid;
output         s_axi_wready;
output [1 : 0] s_axi_bresp;
output         s_axi_bvalid;
input          s_axi_bready;
input  [7 : 0] s_axi_araddr;
input          s_axi_arvalid;
output         s_axi_arready;
output [31: 0] s_axi_rdata;
output [1 : 0] s_axi_rresp;
output         s_axi_rvalid;
input          s_axi_rready;
input [84:0]  mac_cfg_vector;
input         gmii_tx_clken;
output [7:0]  gmii_txd;
output        gmii_tx_en;
output        gmii_tx_er;
input  [7:0]  gmii_rxd;
input         gmii_rx_vld;
input         gmii_rx_er;
input         gmii_col;
input         gmii_crs;
input         mdio_in;
output        mdio_out;
output        mdio_oen;
output        mdio_clk;
input         ptp_timer_format_i    ; 
input  [63:0] tx_1588v2_cmd_i       ;
input  [95:0] tx_system_time_i      ; 
input  [95:0] tx_timestamp_i        ; 
output [95:0] tx_timestamp_o        ;
output [15:0] tx_tagid_o            ;
output        tx_timestamp_valid_o  ;
output        tx_1588v2_cfg_err_o   ;
input  [95:0] rx_phy_timer_i        ;
output [95:0] rx_timestamp_o        ;
output        rx_timestamp_valid_o  ;


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
iGDe174QOvlGg6aywFQXo7uWAhN4/9k0obvYWOWGusqCpX9dMpkOLvV7wn9pURJJ
SVc/k6ZrdDNN54sV3nhuoebBnew1pJT7xrjeSzcFzxk5klM/XPFpyB0LuSobaLEt
AH29AJGazQi9huI94TG7Uid9Arrcpb8c8zYWSAU51rNwORcwx6yzeWBNnYzBaEIW
3Pdv72fMiZwPyCaHLc6l4VLbXh7eqhvCUUDZ6vVDVPZdRmqR04y3M3R8e1LIzaqU
WT1w8/ICWtGI1T1T5KAUprM9gvKBqTlxa/shvKs5Iou0UTuWvWaWHONuz5HY/E/i
WjSC4J10hdZZX/ROXMGQ9g==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
l0h7NRg/On5Dx1GbkkoiNzM4bC+6eT9ViAio4lpYNxma0uN6wih4hhZ6FxApwRvD
/2z+8eIPycdOWy0UQi8jO7G1vIsxHrh/drjoKGuNW/afFzmuH6+W8erpvHj6o1vc
P6gVW6u0emiyfnga4TCrq4yZyriMaa8UdwM5pNVqnog=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
pz7npZw50nuSMdaeJCryzai6+SiicxpMF1Qh+kW4+9sOm2ud1QLskWgZuzOP3Zld
eDRuqoVvyHOrKEnNLe/UOn47reHUx9Yko7viXaJ3jVCCclgNCvPfR1XXCt9SX9pW
TCYnseV/NK2Hc9FTVJXaGNS1uzzpZu38P0xSq4q91NJ610RD/y544HU7C6MVDl2G
ZCMhdFsoCkzX9kbgj+iDM/UVbXpbDQNmBsYjF7MPr4c2LFDBfE4jIGcS+jPPOnbY
O/cTt3YySriwPCkHTrl/pbxcveVfetL15rgrUhbGnmCaiRIoykVRdxAr/DtrmB37
JaEHfnO18/zyeqy0WB9XVw==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
1uCh/WCyGsSf/cIm05faD9XOK4wtO53xOv7TPpCsbJehpJAk+BM2vlto80OkCl+g
30rCL4ZAUisOCxASlNIX1GApgHFDx2eA47XkjmaX6gxjAIw1OFxTfX1MLmEhqZ8a
plbMWGsLxzRQWtzXt6aj0cAlDiHsN0t+w4H/qDZnpCA=
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
mVQwPFmqTyJ2Oii57G06nfEQmH03W2WbdlFr608tBLW3BrwGiZwaHyWMGX6kaUae
Kcc9fIH4x+HLZoFxEf65kWfFxrod45JDOd86Y/vNIq3anZ4smHca5j+E7DtqOfzu
mufzbJLWYC+i8+moWMoXRW9Lx7YtLkO/ne/dy5PEG4M=
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-009"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
m9qcOt5lHUz/F+lrpf6AiPTCWKXE3qqNfJG/HFNRiZ0nckVPx97nc4RMEMTbPAlf
9JGllIgoMFJ7ZH7Ezb7aOPNJkSQm4Bk5XljwMlN4C3xCMI0ALM9VstD55LiHiPF+
RlscFeoorMmSjhfzHHXPzK4LuaUOKjgOInTrRS6PuTI=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 5536)
`pragma protect data_block
cUizKmd7oPh2xiQZDVcoDULaULo/ujZXYxisF4CZzEf3LAfghCSJUPUFDIpm1ysD
AwOpyOVdkwpsbHFBdKLyeHp3/ukdAcLGEZDnW36p50d6Y0AK/dBlEdov+EgG7/pe
BaZqenP5W6M3rNZFaTJNkPkPWBeul3WxihL7+bGa+uSpvZbYudAodr9o2dVbrO1h
y7FrhxuJD4J31Rg/vuDUGXGC/6tw23fBs7xlRLax4NU/eJTOBnQDGY/2jmV39j+w
vRbGlrspjQhFU7AGcQQDwLe5JP5oROtBQ7HjdikSfvJ+75Nm10huXCx6RK5k2wfs
qnBK0DvBRuj270m1kuOd+0PZmv6MCXK3TUT/Vde7PPyBsluigGCqOuTlBX9uHy3y
GBYSgmRCO9+QXhPr2tKcQDe90lSWI5igsXIcFPchS2YO3arEp5GLG9Lvmk35dIy1
O6pp7RrIIVnaxwkWtQw4gDsFhPOl+jX8gOY0f1mTimCIwGHFYpOXP+hngaJlE6w9
kO45jpKBDfn+9zrfJiuj7vpfeo8HaC/Xoivl5ZVGgpwfk1AdATQLkb4YkE7B3wZ1
nmJu6wmUFgMZUr6I1VqydTg3t/YfqWpu2YXzzeoHn7bpKmtsUNCIY79tP+dGZ1BJ
bcX6ROllCP5KEdksQUmKtXVFT5uw8mQx6o/C6aVhRRJqauopdsJcuIDYZM7a5Ihw
oalG5ZFqnPkn2uX0ehbxcxi9LRpbay0BJw3URk728tz4+xQIByGqXUIKMrJjJIJN
Asl/oR7oLNWE/zWUb1nuqJ8YsKhnKlW+hJT9/+uK4JUA6tb75QoRR7Vaakngjywu
SNB/zJXKP/w4l2paF8Zv0pXRKhnr/jGjqC/Ehny6IQBInfP4LL3c1ShjfnvCHWZF
JG4QADT9rjL50Ryd2lJ4qB2gbnufJ+mOHH+IEhF+dCxU+AoTLEkOC4Eo/LJ3Rkhb
REdHsaxfJJPfuMHALbAy2xd68x48HwpA3Fezsv4vdPEkATJ1ktOIPZuCH8+M7coh
XCOoBfflBakhYzAvaFbQUt5IJy9z1EqeLiwuBNyIdcTNo1Dovgee8Bcb5X4WNcP6
wSmfbTuwzNhnKktPjw5WlvT5GVmIbrfC4JQB6Zrx3TFeFjL9HiMg+LS6Y+xnqKVg
vY3YT6SBO21uhc2aap4fRSBJxqDp3WRbydsKKR0QmebdYpC6eYIh2R5pj8xW6JP8
Vy5U6C2Rm1X8gG/5uQ++6gvlealOP+W7jKfvvo3Rind5cnLUIXrPEOPhZEFVLg3V
eemqpFOW/BRkZ2uRQlFlpSkYCsODd7LcdORp3YCB8xFlnqCyD13urrJOtVVQEJ07
apLYpvJciZmsrKW9SicFApiPrkBYSISIA95n0HPjzHHEGkNZfYWaJi8opmeqNFQG
j9PW8AhfiYX6C4t5plreNMp0i27I+VnqMf/WK74HHzn0nZ1fs4h7xWjX2aqFFTU/
KDmt4LQOYIG3B4nuQ6hf+qnwyFTm/yY4J3d+AcnvtcLvCNPy0eEHonEK3OScxfoh
44NxN+hsMBh3QXofCev6x1vWr1pFJi2LEkXPWNKvi9y4olNQ4Th2mv3T+9j/EAyR
PtnPMg95puzsApb5T6KjWiyN8qb+L9LM8quY0eGa4azoBOgwdjCLBWTdQHfl13VK
7Tkn35Yar67fg7EGi6xtyqxA7VqQYvgTl/aRgmfEZsUPEKGa39XHRXD2Vz1x9Zn2
D8GdHEDu6tKH4cauZSoZy5izUGfmoTQ6pme/2I1ZUZPDGLgXmMp1+4REaoqXxksB
KPStcoUA/KdWCEMpSeiwQQODyk2zTQhH8KOSWb+Ciu5ISHSzZeGmcC3Zu3SrKPLf
FCPGE2F9RKCsiepzMa1BHEE8kxeRFqdCpeEl6KlyjWq3U4SRwXzOPHkt9aqemgQM
P6jOuRHBUp1DkRLGjUdI5TW7bVpYNw6xuN+yJwJ43vmBM6mNUkNX3glg9Z/HoRYh
HSRoIzseM7kFUnn8BF+2Tr0sjyxE6XmJH7kBHStQ1YvnieKGSKKbKI8KVGJaEUiy
TENNWKKHQNZ9GA6zSw8QJRerMoLYvOp2YKeoEP3BmcB2DFOU+HHHbbVXIOlQZ+RV
w50AKS0VME38r6K6Q+W9YgnPRQJEEW3j4Ug0/FJTi74AKJ7y5kX6ZUGXaJV0uKwo
s7x6bqhyV9ynOEcdV4xBEmN6Uo6Fk0fkgvxFEhOsXU7zHCzVae1c3Axs4BwIMT9d
QPVDEAq9KUP3882q79DBpKgqv/3SB6vT2G7oOy6RkIj2goNngA4Acd22DyMds90K
ASr9cVuQyHuK0T36y6+4ogJMb+UahVJa8r8Zmq2fqNiWwr1TSgRprNIB3slMEcGp
jOmDuMsoIqocaJm5jD1Bn84JAH5QwyaviYxa77UoDf/vMA+tVp4IZtN6mif7lmf1
aMRR+r8KQbTNEd8BfZJZ3Fhy4xxxQAMSTyncTlMMao6V33V4kc0bE0cWdvHuXzXg
KDCS3/Al7AwQqdqOgoiGR47dVgTgaj95rCE986U+sKdyI+bI76AzyvUV8SQzdcY8
ow+XI5IKKZUjaWm9pH1ODDV4OhV4a3Puc/nWkFUaBFpdly438oAw8ohDODuunk8M
wCNukbxJR8EQJ9H3iLXBtKBC7F+lJ7Rp5j2I52bg/ZnpyYfjGyPIK8prIZJLGhsq
3Kakx7jtZclVeNGf71vCI3QDIxO9Ht6s+wNHOHqjHCzkr9PdhAeGItHJ0uPsNgcx
gbjL6I/LI+vjeYItyJJ8lemuRKEy9fsRI/KzPUQO9vc85zxbcrYr298XVl4mkwez
Y7AZM7AHFqaVyqLfmoxFP/PArrcUnLyLYRsBqiMml5BLHwMywePcY/tX0bmoD0KR
7z/lFbCJmtdom9ljcRb/YWHEMHpfiJSEBZp1TdaCPEZabBITqI6pglp82WZoI5pt
jque/GXIzodxVZN0NpwD8u2rDWlq1pa3bF9SUC7Y4WwUT1UDtUGFajjsOksN3UR8
6VbsTi04VYB+it9OuPKLvl/hNuhEuCVWAk5upcngz3g8bQb2wOjtCNCGjhTKYfI4
n7Q2HvpZk+VEpeUH/sIPeN8Of8iIAvYRpWuj2nLePCJUxXPbEV3iyo/3z4wXNXh0
eYVhc/rZ9bKq5Fy2BK8IxgeuHzU/szWxPgDop7w0qwpxZ27YGyUG09d2NVb+FUyB
bi5h1dIA9Kbqt0+qYhREKbs7mxCu2qu1eZd12XqGwS9010V0f9gC1v2srgnu+f/F
xwUgTW4QIYTbtYBnhgeO6QqFRseSM+KhMYwbGHNygQfN8aYzajleTVY+xg9nRKQg
ZQyn/WLg1Yqfp3jIeqyzoRpUh6Ngu7PGygauD7pmL0TsEAEhhEL8kXZ0hK9t9jeC
OiUZQGUz71APEP1us0WEUHf6YZg5r0MmBD2kTTrGQ45UqJ9ItHA4A2+btm4naR1S
qfP9FQArGy5P5v7dI8bm5mlmAgJ26laL8Kld8V9vxMK/cB7V3t+FFdp7q0jPf/D9
mQYcpH5kjZY1jBFUxJGNNCt8mDYhXRBcj5tgUettiuy6u2C+LYVL2pWMrDJa2JqJ
1Bav9la1MUmscemIdCK8u2vpVn75898zEfMDBEBXIKHkPTMHpuaHFuHiYfu7ZPW4
V43URmyAizX0b0WgpXlbub3nf33hY4FMx+Yd2GwmYK/sEukxNwTll4zeAnadomJT
kGdmB+8RYFxFuPnX4QDzQnYVMXqgjBwgFxz1OQ8jBMmKzSZ2YkDtLCmpICW6pQye
/MRuCvxqC7vmOEvNMgCsKSWAya0M8y1qK/540Q03+s6aD0bp5V7TwfFh+b7TYR0g
cFc2AV8KcH2KXrZVgdzcKg3OnfTxGk9DhXL8uD+wcRU/jtZXma7Om++KqM0iTQRx
EDmJo8hPRC0UJb4y2OQ6OzBSbyNsBkM7PdM/AxjJlwCs5gCBKskZKUe47ziUNCt5
bEeGuU4su2ZTEtVXCZA/3DB6fafPAakGiEK11PM4Pb3AaAdVawJd/l93Hssh2qFi
YBcjy65P0OlzNLeT7/bpY9ZQdDTMofiOzY75XZ/6blqbfPZ/mN2gCpM8dgIOY9JU
wD+yJz+vQG9/TxbVw6owNTfsXI8e1aZUy5HhmqslzInj61pV3VqGVktUgVGIlQLm
op00oU35TxLLxNKfwiNV3+JaPe7I8m0XlQYmQQ+jUciW9Ev6OH+Ds5ZVs2RYSwav
5lLP8Q9F0VHJ8bnLsV3y1OXyFF9yFcaIWGYbm8WkgFoQ+Z+l8JxxXnBkIohSuy1D
dsngSGHvExud3xRyfOWDz0gt26e94lRTfKdUYaoGCPg37Kp6sL7ML9L6Drv2jyxl
3ed43YI7uxUkBk+A2LFZTjXePqxJjXtdrfB+Kgzh2zmYGcU7EV6UPmikhhcCFCD/
SdH+gmSV07/5YtV+QDNVBEQOJFLUwGqV5C2yTQafjRW3OD+LSN31204p5NMtVPbm
mv/2cCgUVt3UQPDIoFJ/NbXtxZHwWgLybvbjSjcNFGSjr+bF8Hxewo2Xo+XDagqm
BZKuikVma5ZuTx/0fjH8THV0cGnr+nBi30JZ4JFOqQkZjXaWfJP624CdcAdtO0Xn
7eLv3Nt8yVQOt6/bW1GkdenQvxoKa9tecL0dGzCwFvuBlvpx5sEcxisWISBX8e2M
L1k9OQH0HLTFL2fOfLvpGQX9u0ztFFpbflyxhm3IUVe2oCcccRfFaB6uQpStpg4Q
/Ln/ARN74851y617z1n9RgjtMdRvxIzi61boaOvuqtpu7djOZTiKRxPY8/T4pEwB
rqouf63O3NopQQOVCe9wg02YZZ/BHHkYpFzgJg7xSkMK80bFZkZLxyTxUzKM0T4o
8as+aoQ62pBS0zZrBXq/8k3Dup04H/3JpjX0bPMaCs5MpyfGtV2U4ItxiOHaEwCP
oVcUsHfKQkKXuG281VgFgxDx8cFlo4Tnipu1IuX1tIef+G6J0UE5XNrkgP/OCL8R
HEjIHCK0BASpVrzU+ViAJD7Blv71NzESs3vy4HL5qHvdUABs8OTkuceP69LIKKdi
04rk7ZEayrY8ImBWphpc8FjqnhG3mHHI55STNGX8grkN9FVbrbMC7F1FXgkSQFGq
Xpn8ZAxxkyY5+03af4NvRNMm/Sh7eQJ2VbPFMz3fRhUY+OxKJ/Ob1qYtV5mZSNVh
7gqe6uEicGq4v0uFLOivZO5eHNbJRZKeAyVtC9lI7aoH1MkWTYEWlcW3nQPbUyT8
23TPQZxdfI6A9++HeUtJyOYhR41ln7K4XNAwGVmbh8+1IVFq42VGkuCLrDqoQHjI
WaYgqcl25D/q+oH4mqKk+SrFgNBbtxJ04jzc/ivVW2TcX0WZH+4z+hsu4rboVnV9
rE0u3dOnzj5pTqmEaRqaYbYOawbFRZynhbCzITQxZ9+I1q8H7WLO8wkwseTpDrPV
g+oBu2SFp7DDx/KJIumaYGHCPpz7dp7TBOSUrkBSQCQKRxWK0Hph/PlkAceqQiix
Pm/SUmHS/9cvi/VhZMqPehv5LIkk5YcfqbK0VpkeSl9GN1BQLxJNhQ8kWjBEBr8+
kDO4EWkRjasDWRoBwOnUmNI/SE0O9gtkI4eWldWPyj1F3F3fdXY+lhrWErlqJcas
xUgH78zcg9MQecBozCUQ5EqAvFV+KThI2fAfAb4XTibxRzT64pXdQPzv4XUMb/Vp
mNQOIT/dGwcuggbWEPEZeW3IRyDPcH9cgXFJnwDXGqEMrIpN5ipquqfKHpjpVpVF
q5zlj0PyF8cqhDKBuHssnfm8IKrh/JOSGBZPHLO/u+ADvF438dz9jLUh4j8i6H8B
0afsa0Ni/6wb4WJG0OlgfKjL5+nygDYGHzTr2v4aH+EtBqAlUGhlOo6QImNenpfD
Zq98yVNSrRQ4UamyT2NlqHNEneAOeq4Emeh5cOSsFpQncG2VSVB2292l7fbqV0QJ
j/HF6VWDU2nNS+5x82FjPIK/EOYq/NM4qAxIzNugj49Rv6R4hEOd4qk9V8htuRtW
Aanki+gyshF61JYmYutIb+eIT0fURxl/GFb09jldYNi57RRSz5SIOwZNMna17HDg
WxUZ8/rr+Q9oWebzD8Uf3L/S9qXOUoLpEwxXvfp5APMX7ToW8/SitkZPIjEHQLF6
JXK8SrQOOKTLrCpbQOhP3KMkzuQuJyLNw8nTbaizhFtYk+y6KkrAJ/qsP82STs0L
OBKZmzz5jUOQIdwUMg9CFQfZxgp40EXzDZoOCk0UxDOytttEAIEjI19Ass3Nqfqb
UoppURwlQ8pw8h1oywqbNm7Uc21+jbUskuhPr26cGI4BHfgPcyB+y1FfoQ66QsrR
fFfgmW7veg47ZH8XTE01tEIHDWvJRuQ1ywbPM5OGtskfKVZ51TL72weemIMQEy6i
Xv4h3IGraETRvmBtsPcIfxk2XQ0a5009zI/FBerkU1dv0ub+8kx2ONyniB9TYTmQ
vE8cOF9MxSAV2r9KFmc8nz4PQABoQrJkFMljEI0ajlQjxPrsSy8udy2In0UXztPj
grdLf25HdTRZ4iIBOvn39rhyTyiVoBWh/Zjt8bDJ4Ox/uJkFzXG+PDmowEFhVfeI
nf7LSunAbSxDT2OxtRxJKmObnkorUYSTvnsrY7istTvU6TJDfgPsKO1FoI0JNUGz
WT4LcgOo/P0RlQDOc+UhfkBWvtE1/UjXnihJFsKn+YpkQqyFziymHh3AeW7dJWUY
0i+EO4jx7p89J7NdetQ0obA808pUyuYPzOiNsSGM8XwVJswsAFpdwzEDYNLRlrI4
vH4Je+yp9gyttTIzyV9FkAMaM2gPLAneH/DRIzh8YQAO7WnuT0BmxatIMSSM6BcE
Orc3i5jvDSmUhX0fbqTh7NEUBUCAEQGlQ3pDnoEW4+ooL0XPe4vLCq/xo+ZkCJ6+
LXGZgkMGE9gRFZEeZ5neHOYMykWmFLBOTY61wC3cDZjnJHWesozVCtD9SHFzAhDg
Zu3jiGHVk4Nqb0rT1qbJ6KxSR+qD9HWpa7qwKzHH+PuvDw09EJzpNNWNRckmnx2N
TqGGBfu5R75hSqS6PfSWMhQd9EkvmBE0P9EEK2ib0R1t3hgJoVQFpnCUz6TW2auv
a41ykYBhWGvG5HBqW07zoFHAfpIu2j0JZRfOdzdWPRwuTWS7/HJAG3sZNzpnUWvV
jCBhdDH4cYhwMMgR24Tv9Y2hL2vQI48a9pAP369re6gtyQAHnMwot3iSF0j47qza
cGY1BdGkg677rIDPZ5MUDLshUy1H8+C/2cDDSk01zba31LxnRl4FR9mJNin3kZxM
ZzPGoQF/RrJB8nBGgE1T47J09fTE3paePeFhWoeCHKviodRLar4ffXcg9rD1QlVh
qRwBvR7zkzxZidJtGixRxQ==
`pragma protect end_protected 
endmodule

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
cbmGg1yiqOzlZTbVYXLPLT6/vDNIzKdVp+cAXtzKATDo1qqPwsZZwW0K08GnpHNT
kqMSXqNu+ko28KGe4/sz6sbJLpYb1A6KUDaUqNaPRdXjm7sM1Q2m5/bp+ofaSRuP
03CfrVX3boFCUrS1MO1nGE7YgIAuJ0aS5G/9looGyoDqhd3rv7ZSD7+sd9SQwj/V
RaJLHt9uMopUhuQSZXdEfyfZYrAIEZO2XOhN4XnqJxyF+nDEkRAGujDfuBijoPK9
ndy0ADQfU1qYjlUKaNypJm4GToUJPFmGyVC+w0x8cu6r384kBquCmQIzXjGkiBi/
D3298voH7toy5EheRhvEFQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
nW6+ihVzfoQpkFBxnXVeI3eCD3Zf6aPpmhrYGTMke41MAVrlnF7NGDBrYKpve7KS
joaaLg304yBlr09It1MVsa7x5hoR+uyXGuznPhvKsKs920QmYkw9XR31Q3l61IkG
ENFp43G+bt1/Lj+IkhdYaMsFaL9IYyVCZalxXxTFwUw=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
jMtncoOPZjlDBa3wOTne2zFc/eA404LlfePFlVdDanf/Z2v41z2uC8I6vkKXZyUE
sousX13rzpKZs95eVCpg0825NInD9jgSE/Qiai5AVd6EHqLSIUDKZIfiq5pIomHU
1T72YQWjG6+KPCeAueG1hDEKjoYADAQwcxwdolvg8FfrckdEGXB7XWCxq1MJskBt
MoDoG3N2Chxe8Pt9JXl7cBZ4m8WHoTjeGLyZOTbyJHdiymQmNCwPyN7jLYKpD9W5
CBsOkgU6jJK5hyn5J3QAo8qCje1v1nfbE9TsMTXI7jFmQ1zHfvytLEkdCUWTWFcS
HSqp8sHKKj30XMVrAv1feg==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
OhQd+7NF8cE4fURNw7fw2gP4AWDM+qQSoVhcOAnAdx1/QB7Pc+dqhQS2F94V/ti7
itnBXE+V4HrJrj/E6IHniVakgJylxk8gRjYR/ZexcOodwyvW4SKWgsD53ELjn4W6
YQXNAIuZWIZ1yD0nGC9rVu8uz1gAV0hd0L0zwvfG0wI=
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
b9eIw/SMKFlbEJElLAm4haEyMwMVKrauek7KT1OLGSskrfKqUk5Gr6l42EnuTs96
eXyv0tW4fh4i7pUbsegsjfZCnq2KwLlrq86LTOS5QI87+JbvIDc+gwdSlKNZF7W3
2Vyc9rp9Mpnt1pVrqxHBtSHofNO783bfyM5WSquMRMM=
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-009"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
NxqCKW1wKktQG0pPnXpNk3F8TFS1rfXsqQS56eWnGTZboT3wwT0wSEuDA6meLi1K
TSh/bCGcehADrWZpf+hwpYL6EPwspsEywCAylg+neM4GzPZPrQCA0K2FB57ZVsTV
29FI2jbBr3ajpp+zSikXSfFDX5Sux3n9qdRNm4MsIdQ=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 325280)
`pragma protect data_block
9wGI/m8Mx0B52Bsr/lOho1RivjyW6rcf41jLUn154A3UEI/IyVWhKe/Pt1t7phhr
obM154YSrSicJrvy2EeaKkuXUo1zU70QcK7N41CvUSLJxvh1MImaAqpF6pnCZp1E
K1vnE4SyLtTjwypTrvaASEs4nGiT0+ZeViCNTM7q/DxCbanPnfuxY+ChjT8XtY2l
1KARgBy+7BgZw3fXPJfAKZdHmiT9ps5jpYjDgA0NZP+VLOeH8mpOGnmSOHmk2oFq
BLBmHD0NbVecytyTB8rhcAycdDiZZEUK+UJUQidplJ/w+XHiVjYbLnJul9mMGttu
1Tjrhm63RsflCdnYIjrEfvny5qJP1eQ/8nwxHpsBm+UrFDoWdV2ALnyEV+JIRALi
lX7D3cjnxoJsEMJ41hpSoaAawB/vqw5a2mVLnAlBI66Sn12ksBKvrGkhe9oEHi1E
TyNs2rXm29k2SuZkAfvNf20nrHBdm7XEdarqMx7Iwuo/MytJLH1oj9jqjm09r8Mg
wMLri1Onp2xWDjLJKhuIsmPSGW41WNAbcun1GjjGpjAIewKYb7BbQquF2I/z7+i+
5KOcP/XwQZPULHIBygI0oR+gkWfHtPrtqjhUMyfOvuF6lvJNTg4yTidFlYNCxOaJ
HQW5plA3XyB9l8xI4UaVncaAZTiS5yUCID8RkNHeg9LtUmler11p6qDJxwDhizgQ
L6TN0U1A8g4CDS3sBO7UsbguWXA5WIPfNDS5E/YmEZuR+p0VASdB4psJROiTBzrX
VPJIL+vMJKuuUvy/0+R4dfzmFDt62jGxvHC5bEruZa2uS5BTFKR6EsWjW6+D/Kcy
Dh93m590qC1W6FvnxE0SArgPn9xCAPXk4REcw7aSN/PVHz61SEMnL7jlvggLL+iB
90Kpa3gv03C014EEGFRs4J8760NmO4+0MQrVqfVgBarkSOJVOLnocbg/jSzL2Jya
pd8E1NpXtKAt2y8EkAT/G7HDeQcyCji81pPMF22BordEgrbidVHTgfekMY95id5Y
q2sIS+c3r23gb5rHDXjTaBAc1uT3aUlyEZWV6vwZu77H+urlCM5Jbm2xamuzoGVu
AHJzTL5CUHQD3gjesOa34p9x/ae+UuuHl4og+BVIKQ4e8zqLYAMswZTN/PHTNsuY
QH7yRRs8KJpYP9VlMOh6NOTdliE4gYbwC/U0ZOf5OTB+MjcTacUI+PEAmBc+HwwH
adQMppWMosJG4mzZQ3TLndOB38FMcInsV4Y3eWn5JbT52byqPQe5+H/trc69ED23
5/fXPRp/p9+gI3H1qbvaVMQBpBowcC59fKcPOQQmPr5Dr9UvT1J6dI5f3QirvUau
7RzEeDyxgI2Gk5ZNi2k7efjgevHrXccoy2BOuUWwJ0cBmcJ5lGNwyX0ITt2GgCdB
+SQdSqxu1yMIBR2Yf+x2qTwRj5lMzRpzC3zSMVIS38drDtbDRp30QJMFMwUSWabK
D9Csim/qNAbRlJi5+mSIa8MCcw9vFu8wFPG/3DGbYFLpxgpfJudtRsDy/42KsclV
VwoKOg/ML3Xz88nP/A+7oCkUXkiLfYcTYDUedwsDwhQ28XVU7R0+PWjzRt7d2KKB
9Htl3oYlgFySU8cE54caQAyC5fz4x73saByd9a37JNq24zm5vAfdp481W06VGF8D
WHBugMe/AZNNh6XpzlEdDbo0MjhX5NcownkE/VDZsTyKOGmHblCDVUK3rXKfKLgc
V5O2VZjV/Ud5eTKLd52+/QzYl8F+YJJ2nmrzRoQqzoWLhj+Ug4TlB/4s4cH7Hl3+
1HugDuwvHO1RRG5aOzg5r7Pi79F48G+kuHonReyyDeeboM7raaMktvj7p9kAdO4y
o+1BOHl+n2roeyL4966oZH07lGYK52Qognx4wiEyCDB3qXlv0WK4jF8Khk1X1Cgm
VJx3mO6uzRJcsJoVcD6oRQKM5EGzeZW0Y1h4RQbkxq4cqsqkGCcCpaS41FA+hOy/
/+Nr4wGEFRLSf67USt8RsV1/hCpwlPdnkWHbOjmycq8V5l/7EsD3iFd64PCyzZF0
LjTo2AVJSd0l0aXI+jknbfyy89n8FdvXT53LJa8rw3+qOmQx0y4kD1Pr/X1IXGcJ
DdHpE5caIO21BVUaGUNdLVcp/E6W+kr0KC2dn7lEp9Fh1uDtPcLvgI+Av8iFBmTK
QSJ0jX4U+ECOz1Km1QlwMt6E7WMgCqkwpJZGk1OCZKbqmWmWHaRiMA/EQBMx3OwQ
YodaouJ3yXqblYFfvhh6PuogWdXtDjkIDW2OP3Osh1O+kMMJmgKPzhAcWA5Qbv+K
DeqyJxwJvGnCDfOjQvRLq3cAqDgXQsqIr8xwcuJG56Wjdvzh4rEM0Zwf68BucKMa
/X9ycNhGL+ja/FKAn5Gbvnf5UXdHoSUkA/XlA7yq8CdpU0V+QbkXUjUSpdD45T62
EHMxEMXPzgvg2NsaTAmqG3mRIUrTRzwHShoaCFzuv43Y6LQgcC7CdbbmVeH1kLiv
35+CVUuwB/7LuJcxNpRQvzflIBjjFhGMZbu8pAicaWxUEKPyBrDEkxBohNvQoeKQ
q92pjQvyBHX4gY6GE5xwmwIQE8T5KpxpIBXsccbl3Q03k2/E/dPU6szsQoQubCxl
cXDuJlZYSYTVb6aaRVixk7BuYLyxOsMGOXhwrmZjzz8qJLDuPKpHfskHzAlC0ojK
/7KDFWH5jGhvBlVjYms583FLtuRVzX3xih2kLs6+nt75+fps0cMRORClVi/qBbwO
Q1pgvHt132nvj8BrI9KzoBzJgMnNgr/zigjzgFoqfiIlLm3r4A7H6PEyhtXqBuiL
QJmFPTyba/uuemkyEaOu4IOv2tAE5+pe1vdSOjjggAQBpYSbn/0bzFdxjgwLMsmM
aOXPF6InORTCAY5kOve8Ml6luFNrXoUeEdRE4dVPA6/3gjgBx+q7ILSn9vr18P2f
WxAYwhgD4FL/NvsAe21Krn0gj+uFJmdTQ66cZvAsVv52OXieq2j9OY1Mbfb24D9E
d1JSsAWFujy9NLkqLU/2gUqBiCdiO0vlmQ9WJbuDblJlqmOm5hCjFJu01ZEPxMKY
UEpNqUKhzy3F5J8cchSiqoszujkOEOp4/FGkL1xBW8T1gGqs1N8t6h4yI4DmJF4i
A2CEiKHn7+QDPENMuVIB0MzdQ52U8Ts8ZBh2jjpFHin/EwmsphS6eU6zCnn6oPaf
0btlgBo7NPlDp/DLDl8hMTdbHsj0haixDmCRd3w5TEhB8an2OVHDgCcvMZascajw
P6W+ZEz1OUHyZ9NQRkggZW42GA9bcugwmQuBCPOCY+snVs0iE89+Oi7ac3xLF3eh
U7+yfEKQwT4tpb4Jov4+QXLKI/yDqieyWw1qENjGxa223GKJkRUqTUmGAqEP8V5t
V2CKjgIasY/szlW5ZGd15vPGFUKvqhzhM66YZeBM2KOxwQ8lC+sV+7aTfQtxKP16
ObRR1D/eE7b6dHp0chRJZqod6PcT39xhj+SNWmUEMdMMH4neXUXClfgejXZKPvrS
KxGeV9GxdD+u1W0jowpcMdVXJqy85D6KMvRY42f6dErG4G2dNN8yt/c8Pmo121xV
JYVf8wDCCSlKeTbKsRQJ5DSl/CHau36ry1tfgcuKFY+goRYwLN1BQeiXmWCX12f5
7jBgvxzQI/rPyl2NVgp60e8QpzRdQoOH+IjMkRrlFW2rFx+I6tpyjHgBNrORgJRP
yDy04lsINo2CwrDJ5WjpdXSyx+Y7qTN1FuKykFCjOJINgjuQS3eyvahMbMWg7hIR
TnCOrVikIn4XreNpEjUefCAQYggAgJCMhJ+HEcTjdSsnfHxA6oMvVzxo03G5s3rL
ETHEZyp3fXnQjdtACTdZfgA3nn3McJ30ePsdLvrVVxt+YJTc769ZqmvI/JzpOU3Y
s2l1s7HQtAxAO+yEyX4BP0gfZA4lnaGxIfh7L72Z5foLj1Cik0a10Uvr+HV95S5n
DTj95vydC+WMIlt9gVWdAp1FhXqHLIt5j48ZhYo67NiwTVsgJd0FQ9wtXSr4y3jm
ZcO7c38uZBiqIFfT2XRljAG9jE4v9/7IocuFD0RsN6sl0/uRzhoJe+TujeI4B2+c
7PxwsIZIztb91MmAQHF/kZeM36AIve4HPKyExfqRlb2t7Z+kgR6gbCkEAEcpNw1l
MOINtO5Vq/OcenIdBMG1ETHXVyBtsP9+aOJKuu1zrA3LiMtR/R/3bVhDSigk9yMh
/INnFLrulwt06Z17JE/C8EwA8QEMcjUv4m9OqiIOo6OmT8x8LEXNmEW7e1/uzba6
Z9qfaFsNBoFhFUsSMdS5iJ6lto0xQRyjqboqMDMBDJK0ggmPJhaTzw5UqKC/cuOS
WwGZvianOMWYBRq+8ZkKK7PHQmbM+K15eV+NPZ7JMbK2eImF0q8C4KLxPCrS1cCq
efCiCgrfvtez6M9KPTSBANm5X/XhRGXNXymWX33CSptyI7duobMA+VPfwnVi/fxS
EYPAH1wqXe6WJJx5zc+6v+hj5VdsfoYM1MKIuMo9c0d11eB1dDMjUSfk4Sdg7EgT
U5PZFmyAGponJ54gAAJNbIRFIW3BUEAiUcEn07bQGOzKbgMnlXNGnnJBzZo5qc+b
Bh8FlpdjGqSbm9946tNb2bWwQYTN4k2wdMMwNnhQ+VE1F5Kw3fTaNsIiyAWmOMub
JdUfUkfxXugDzBrfQ6ZptPymEfeaRb3kaz6HImtL6SxzthgKyHwR6yrxhL/D8tLi
H1WzgbKLHTduWV5qMKrf1uugb9rcPYw21F+2cVzFamYGt6mFchii0vEMfWbVatIj
8U7KWO0OamOWbn7g1ua7I4Gsp/H2s4KB3zkiHaYrYvbzJiyUdLBOYpEQHRqKKpfY
dV5+zvEWS0ilvXnxy39Lt7FBVhnfdlb8DP3Ikd961o4BzZvdDkQMnF2rGgXZrmtY
Us1EK5xm29x7mBCGK6U5uw2qLpkHkTfZ32hdqCa0J48jOuKcURenrWMOGNBmC7e2
dqdAB9paDjPh0pOpL2B/YRUVDayOLVsqw8feDPEuCsSfsc4gKVbKqN0SuXYJRSvU
HPSIl7N2htleDuplrh7bT3Qo1oUYBovVG8Qn+uqVb/Y3kewN9rIi2g4Y6RWCuwE6
tiCNBUdVk3zL0XzAt1Ze5awhppCfJECB/jWMvT01FrvQhUGQCUUSJPB838eC1KeG
RQoYJz06WvoJ7jb4SqbYwtRo5nblXHDrXOa0lDbgpmX2ksDtAG1oS0d0wIP1VnP0
xJa17JAI+KdiFqHuX/HDFAvyrVkb/quyG4Sct+u5yFFXjH6fvTGvAeJfpKkXu+bP
ZcB62Njv58C1QKPwgBN8yOMtEeF0s7YlA+RSjMv3j83ycLNgVwyXERILvwmp6vz9
6BijCj9h3EPU5CsaJrEOv2Qd6glFkntTHwk3eFAF5tRMJKpOZRKMITxRtgVM+FRP
plfzdLZUx3SkEevp5EJYb3Sk4anmvyQUzy2eSvKn9yHIDwOQRIm5UV1W+7eHg89k
NkU7aub49Fqejj5yta3QPsk/Jj3IHzVRiEVxNx8oNop/gTN6Ug6JfkqJCCakhFcP
e6WCeUBhjyU5IeDiHhA+ED2uZrhi7AxB/kx+PlAMkkzbu6Foib5+ePEVQEED4NTT
QNEDsu0su1PDMjqEA7Rn1pbYeKFQKrESzJGGGh9zDRM3vp7Wztu/59uD4ea6OR29
fxAu4A2tv/ny3aGIGH2L9TE6vshLe6Xhkub9HQ/VdnzuIqmSlOXNiADmerDjBnDi
udckIR3JLAdNue/j13LlRHSp82ccIL4luUcOrjeE9zeGvo3Zc++qj5rMnC1rTdGO
TXWZGS0JISLb5KvpQHCxb9tt9nQF9Pek4rAjdTwXvK7tb9iKdIJfcm0F8E8fu6Qn
nR4rPChhsWY4TuxCf5xZ729nDwh3Psz/EnlRvTsyzzu2u47HXPROVU+JMVa6b3XM
UXPx9VQlUEZIk705nyift1xMZ9E7zdRTFdRk0nQGLWnOjrhpR9TpyZq0RvHK4jd/
shm6dWM+vckewIPlgu4JtN9HKyN5wp18CP/N9mTbV+FiLdvhwUtiBo71rx8p0IFi
2Y0+NZwuRj7XnXIfkOEcJX+ZCJOLr8qnn64uZqmx+VLtriNBRs3zaBr1Schpxalh
CHK/El1DX9abj3bysnB10aoN2DCbR+fPkvO1BdYrK61UoBh8r5KlkrYvibQCH6iw
XA9blAnZNJWWl/9H6aFW2kGHyoAuF6H9jZBSOyAwRbnswx/rWO3pI3JLpwJK08km
ntjfhbrjILh8bksSBNN4TmtQOFi4o5Kx+qBi+AOHUlFbVzISTbSsEU24zrO0Betv
8RqLtfxQjAurjs43uq8S0ADuwGwtpRIusvff3VMEux7O15wO4d6iauq1WV0b1vdF
2jAoLI8X8/cJGZ3Yj5XSKKuCImMESQKYza7vCUMEGApON8y5F/5BssBGnDMkdzBQ
bTK4seInqWL4bPmxi6vfdkTYvOT6HeKSbYlxH5J1y8qFzE751yElLrbf5Jj4Eklb
+A4wNh6j1W5jmxxxky+ZpHRU6G15JljVe4I1QoMDZ1+9Q4P0pgbRW73OiJCHQC8N
30ccWWxPaKE3Yzjv3QGdy+jEKJ9Iq489kzA2i50uZEHW8ZDRz0R4Xje0xqS3+fBQ
V8YastHz3Aje6VxxFqAaOYKPzxmPcQOQa6oN9YHft3c5ArqG5IjZQlipUno/288y
+VMguXhNQjKzgwW+hBNWZn+/hIkDs05IBjaLnrMn39Ogvw18/iHL6nDWTUKqidd0
UNZ/Wk5n1eWy78YrvomPpQoF+g7UPA2J3TDK9peQhFwVXdtWuD3cSJmQ9lp7kMRr
W4Ps7XedOv0Mv7zip7QfvWHdB6QzRkizu41IPSUzSNgrbZVtVyo5kYq/fcWZZY+a
qlEMQUd0rU2pmRwvDMXGFN6yKs7TMR7TI3+EnuZgEucaYid4TN1JesGG1Ed74wr8
fVU6QnGtQ9ITV8sDrsGYqZWb3twt866XuIoRW5p98/65rGySxbQWVvsAhPgOREgj
gxq6rEYi3ZY3XEM2Mz8UX9zFhQ4D+X8sPmOhSR5jRu24xepUnA7VmspJvIIqoznC
FcntceXNPSLDvdsln+o/72gndNkTn+WyvIcHqXXKw3uftdSRU8LCJJXsdj2cMWIq
iyKY030y/LHi63hAr9H43xK/2IsJHZgQ0YxbZj0lHebBO7tNraECiQg7WQG9bDLU
6ezT+rZtvVCBcpAJIS6opDXoJk9Mh3H2nOX+1FZUenoBurflinLGB3HQz2B0TO6f
b5rz+DvGPFHjOhmGx1lozxUzHCjKNczhKr4B/9sEFidarPJqGT1Qg6XidwKLxmwR
5WCjUWpqVLGyzJVb+qDpV9SqR1bnHptypwBCXt26+dE8orJGAInck+hzsixiuK7D
rI/08eHuaPT0F5fcoeGeRpHLy6nyEvuYpnfFRmvfi5X6b/nWWZKDJ8GNVPq9CRC1
P6wSUPQ08PuQeER4aV/LkxGJ4V1GM577waAp7wBQKxCqi9sLERrexALzKa2JfRQ2
QMQu7vTJ/IgmTKfZrrc4GuLy9tWS7vF7XnEKepv2ggS9tftv4hu6IVLA8SRg4e6j
viFeR/59au9WKKqV4Y6FNMfIYw+gA4P8OtKLSxtv55DzFKPpLtFw9kC+OB4AUbny
zIfJ021aFWxF+ck/uLJRNwjv1CiIwW6SFRFuo4ht0G89d5IJnhvPvrvE3HceQ/s+
Tq6pHohzeuvXkgGhVIK9LLYflyTkBOhuJQsDhclv09lCxE78EKht2oOspOaWFBi6
oelCVmsi1AuaAM95HNcbtO+Kmqa+HZ6cvsSMnu3mv+xxgDVHOwBMTRf/Bwxrie64
95e2zuE91caHmKvXvE2BJtv+gJLNKIeJeaLvH5uGT9QEs4TYV/x5lm7p64uWT2mQ
PUqzLSuaYuYAOQj0dUUpIHFG3L38AaSNFDuyhIZ0HTwUaN9bkapBw6Eqm7bmV3x4
PTkgGaN2HW58j4CXuuqaNKlt1xOUV8PPC2qVPfU6VFFiTOg8qNeyYUUDUw3siLZG
XdlE3MuOLDdQK/AD7i3jtIAV0ToUS9+FrbKHRO6zr/Bf3YuDcGbyuS4zeNI3oJEN
cwVecBogOA8Hsy8x4Ihr1821fTQYV28/+fz5ttRWo0rtxNRVA4+IUx2uafqUSQcg
E/9DI69YU0OIeWtpi1FLxUJBsJqihfLrOxCDc+fp8l6MkH9efK/hybKOBqC/OUej
2Mdn2+GLK7UmkN68yGyUQRjituPnXxB9PCxM4xGzOdd5cFys9lmV5Svnj80lGlMs
bI79uQf+eKqnGq6kOju3wYEyheVCK3xQqCqo7VbugbIbCSCv980c/bo4ueU0tWrt
Gs4kDBt8p1nH5RcsA9vocIUWJuACvjoQEoG+FNQVwXbuiXi6rPihg+nGrMsbVjSl
GkvXfbx6uDpCnTmfgzSl2ORsqJcjh8ti+IqwQ1evx8fONGuym/ggjJNm0LYAHpbq
OD1FiUj38586CpqVcfLO41nm1jsrvboUZl3nEojEWnZyxX43k7KgLoaqgVYkRCB4
Xa1bK0INfrQtLPfnMLdmbXKbCuuB7D+8yolOij3T+MtuWRtv7apf0XHyhDR8Dzr2
bwWERkPsz7jaGBtOmd/RbU249ElDw6TLbdRYPg1bSUVvTR+D+BlwlNLfh9lPoGgx
aU3HDHETD6rUagb4ZkwIZr2PEkSbRHiy+am1Yx6rNHpfVxV3VgU6wSCQD1E3MK5u
m67YlfdDLVsQit1ntkFBpX7mMh8mDNGU9McVuk+MguW04o3+li1Nk+Y4J3P4Aktk
WQSfnWWtYXN/c0IVaaFXEN12bu10rIJ+LCKJ6/qTeBX/hzTKt6RuDo6PzrWd0H7P
Htnuoq0JzpD/GWfpZvtrZeAD63n5octESFqm78eccJXtB2P8ubiZHeAqwFFo1BJL
gdUm7InXAY0ow2wJmM9YL5reFbkHaB9rKqcTb3FLjJRmVXaXdXOhvGH9zZ4Mn8mb
xtAQjxtCklvfRJFXXBnWhFLSDSI2T7r8CIozyzW+Pk+ekDC08flutuLVM/O+Vs1a
Wt+pwKmP5FnGp2+UIYOlEAoqetdNN1kCwKCLcd4tQg8BYFWadCU4K2MS2ZVyFJ22
YUVkvDraUk1jsF8mNL9X5xZdg39DNL5bdeCRdvZi/6fg79zasXoLAfrOKK6v8Md3
p88NDWFO2DunZY56B8asm0144F6JZPhAOO3fvzxIBhYYP2P2Vpv1rtXBLTptkpe7
jO/kpEbRy1bB1gD0GkAIp3bK9ypY5x2y+LKh4L0vp74RKwlY8wpZRN+3E5O4Y1Z3
W4ZpjrzQaDJ/NUobIimbMPc52MmpgUfH7qVTGy8jQqVC2DJ+l40kQRhJe9zdpb4l
EaX6/LyolG6by7TOmdafL4bHZAzROA5WCQN7OLOa4U3PqnKE1RF6mcga8xDs3/5S
6Btduyx+iznXlhn+JMKG/2HGEboCsI+qaNFa9liHweaQs5aY8fgxGmEq+o4ZeI8N
14xTW83w6LKxCCqQlrbmw5KACvhPLc/LDlTvCQvNLbsofCq20eM5jmewgBMDnog6
qF0b6qm/Ds9z6a/ieJoBhWfjDmIw45bF/zTJYtSrhMDuQNO2KmYkHdtS8RA7f9xo
MMhzPpIJKd/BJALViNRzVFWQCTortWOZ9bCf0ju3iIpYc2ZcnlzbrSjruJVzpXyJ
73JSsINfB2ARf52Ub8iBpQy1XGTzjmrq1uh3L84zdRdEetMzj0cmU8HUllofCJGO
1LEZYFyYUHVgILFlhj8vpoPnUb2G/WX9pJcwTx7tha26ZDRNsyEQVC6SLg4faz3P
5DRd0rWu9JQYkf3fazi1dl1HcWieEeI/2qCpDg3OvVNNboEyWPWLIrhaQmqtgFCl
/2RER93YAvudpvV4fteaO4GVlGeqz29sAYNXShNYZM859uLANupApZJmUHKfXOOo
r9XLRqR0GdWr0Q7PrNg4IPmfi7DkgATGh2h+8Crzdx+05Qg9D8aMdNOflgvgsWqP
YLP8cZ91VxB0oafrnV8HEzYFZm6inrE4BVfdspPgbeKs6MJl/LZar+6/1RbhSp2j
tU8L0SoZPDtEXXLtNLtQk55sXXNFw1+8bP09AYUSeETkA7MT8Se9YGe6qPGXWkmt
shKifqwuw2yuZFMeOfA3hB6hk3sb/+m1geqxLHzY8TP5wkBu0ipGrqvk+RPWjbOK
FC4CDVCQGldhOChye+EaddLU6ucennOOt56yMn68wiwTKVfpO+CBkkVpj7jKhWsq
yRF19OOg+Fa8SdOwoyYa1hzvqW2V1HYR+UJqJpnJfMH7lB3MgQP5/1OBrxvtnNip
Cap6/jLnHDhXoeE2yGZcmJuR5IFYWj0sSMqf0wz4SC7p8yEk8rAuVM8uMrvrlKS4
Ha37Gq4zT50K0vvf0rNRWxZTQAdon4PzIz9588seaMevdshRUmmoLBUg+DIvQHkg
s1lURH6kU2xU9urSRjaqC1Ti92KlqvF4DbiUmnX1vd6BcxZdHDpkGRbBu+BRJuli
pEhhZmAjNHxX64eKLHH9I25wk3+MkaGbAZftyct7srqzlIqiKUeO697Q9wCJXHfK
ajbjI+J6iPlFJBGIiUT+UixAenyKuopBiJannek189v6WhzmRKXqfmyhPQBJWYVx
NKZ+QgPKVjI/kzvxKvQspnC1Fs3qp7OvCEo15kMJyiAijeO91No93tgQQOGs6Kzu
Phm6Ya1xte/DJqQ5N2UFCxFyDGTWsA9zC2OrZmFD/SsKidjPsce2g+h+CAfCfXye
7j2IMZO+JSaneYkKr9mdypt8r+CigJt/IP/Ur5pq5jCubVEt67OKWTOaSx/h5r3o
UfYVtQbgMvxwTl2YrRbfy1Rdi4c4pnpPoa4yr3eVxU3okWay4KjlOVj3MdLnbyrF
6PR5JaskhxNwYbfDOQuvYcmfYYmc6igRlkWfxz3aFsRYjQkNrJ4GmWkQhgQjQniC
0vNXT17m0z7LXx3F8Tzd3fRR1Pu6q0K5ptVpMi2xfBQ2h656OIBCY80ZMQWE2QwT
fo86SFyn1lGO3SWO4uLX4SR2GHyTudy1yYracOZJYxDgFUsru7Q0qmijhBl/kwup
cm9RUb+PPlWzykdymnBOgtCTR8MZcJNwFwb7+RVQpF1GPcf/c3BoFVT2sfICz6ff
4Z0ID026QfGkeMd/QA4lQcmOnI3MnXxbI2+FsaZpMh7yRsyBqjqGY0/ivPrWbb0N
+9HzsF+GBD74bGsJJ6YbBPO4nTABfgQ1XXp46WqyUGcvfxPZQb+aZQX/47Mt0Vyi
xO9EvD0XF3idtfkmMdg8a0oYvggxFDs4zWAskGmzzrbniUXU3yHvqJz116pFqD6q
7skUmx7FxqFo5OZIq5cTqR+MoN7nj5G8BCtqkrt047A+dnJDscvfhyZp5fkgos+v
8IzceqAyHjgDbgYiJKvPavakv+NrUhpa6oc27jRprHDKTeIWwqdAhtPgMb3RNOHO
hbWOYzzY/wFQCy97mNDsN4v0NXhDEBV63MEjZZkaLSYzo7ypgB+O1PQANUBvb0Tj
V1wh9mEU1KrC5vWji+cPVyCv5JSvODMfcMsdDcmRqy2evFe3Qr0M1FJ6JxXgcMJv
jyH/RWJfK4na61RvfxAoCmZqQmRJM2dtG9yVlR+bCdYhhaw9ewWvW/rh3fYIEpNN
PxSsR+01lGePYdYwpm1gbxZyf2EI07+JZJKmMl2WXP18gNgN8/Vu+hCT4N9/UtY6
429z0wYLDovXnJ58dogWDa22k1ROqDdswiV3prK4XEGfYZYJftiFaL8VcnqNK8io
MSrgPcaGMlrYFxfxAB2rUWxvk2BCBAXKqRM2P7HpGLw0Ga4E/NZgGSd8b22hwv9O
irMLAmOaBdbqUcn23b1OjoKH5daycyNzy+s2yOaXQ4EwIzTkxFHg7z95XSRDOLo+
yLqNXdt9SiKt0wdCZ7gXyNA4gUd7mBOfL5qWx3RRknQbrjuxw3zdo2PsQNnU5Yes
5twsGrZtF0Xg0zElFHarsljIHcLm8XwMPpRTNWZ/qsSI+TTTc3+bLK7ttdWteC6F
hllMZLyuZNg9PAkrxiz01wlt5+kiUcVRa4ZCEhOlDlYF2rcckPT0yQB7HagAM9Js
C270teyn6nZKuTXjPkkvcBuboVelqlEkVega1J/CjtID4FYwgawJpRTPis61sSJ3
SDBAaQWxeTWGwOXHXUIDGD04N2W2BAdwiYMzS8/kVSAfdWxVSyiCEfBXMNIDheqO
29DFDy+QwNf047WbjyJn0dnQNt9Xmyky4+0fbTt2988SmrEJubrsb4xbP7aFCjNB
w2usDOjOOtrQAdzH2sgmq+AE/17hzBF7NiQak+b1ekL9UBdrDBtkTA7Ix5BlRgD+
9ZylL8QMVJOK+b3/VdRtvpYGXAQ2gmga9OMoBl8CxiI3EmnqTqy850Tl+Nd/Z9aD
TK9tbkXKc6arz6C8hHBmqaYwuh2LNIqPzCgma3fA+LyJ1C68fpYdpFK35ZL/RAHs
V/Amhza3OVtn4FCdOpA8952dd7pUX91iNrS99MEnJzeA5lGuD9mB8IQN921pZ4u2
vICzb+zaGtHP1InN3cDSuE+7ZkCaWJX1gC8Yc2JqiIz3uheviYnz767LllUc7QeP
nt9vMmtLwL2Rz7BJbaOGQOjLEq4JB2TVS8q1zEOoqsaKIJmKqTNZRULS/tc6Ora8
vcLClkTvO+PKeOVHpjd86tl2PQSRC/+K6TIvsty5K0sYWitf4QvxoZ/FdFDA9TKE
yR9Kc5mRJx1IEiRN1HkYnvkswIbRRSB+qNZVKA3etvx0gfs1DiJVHuKvRGZn2Jdq
7RGF61cEochtxSFY4D8nDTZwOUT8CrOBGXRT7eat2mUfmHtkWkd/gl6CwIMTAlvg
chqXIyhYpCp123KDwJzelV6sOBY6sgQ9bntB0a9S19xo7wLVd43an2xaVE/hYdS3
kWOLguINY8e6t0HkRwY00Ap2vYjyzDhI0Q1i0bklFObPj4O3ya9iN/6TtTIy13ob
/sclMWCCTZ3PtpJrHb+bULuD/RV8KNSpF/6yaqU2tqYAs5BTyJLPszmUj/vGd7fM
Eju133S6Ga0BBv+JPM76x/QLH79Izio8kVebsGUPuo2Xkn6qyI2X+hrig1qI6AWY
g4PbwuGRGuEmhT6yVoxD/wQtrodu5IaD9y3U+0SPFR8B9FpFpGNve6cuvtgqAfU0
/rG8jnUn8tixev5Acqazqp0VP/8mHFG84MIm4pAeWxYx3cqUysbxpvO0+MdIDsU5
Xe6jTxrRyYb0w7iFzegSsL6zytIMS9JJSvktkbnrixF9QiX3R4pUta7ijjep/6dn
sYaD2SJoldz3/pXP1RLXJc//I30aUqFTMmwzVYY5LJiXvpKDEdcIhxydcadyU6qn
GhnIV/nTrZCifa92IoGGixGsGhUjB8kN0maesayruzDA0+jvfTrqvmWSAVsc4IBX
bxSVNbYjV2r/LKmOhs4z1kRI+cambsRnZS+S4DjmlAZwgeywciJJeYo5sdbGy0eH
23XbvVzsz17SL67ASDGgM6ZMr/UtzxXHV3TPnxWQzj3o9xTAtiY/HpLUK6IuPnrq
BcRaHWyq3R/mTNTMtZ2Ht+dH6U9CZdJObqTQKiuylu1sZRUKMXnzOP8SPAfHlp0m
lnfWcffe8WPhS23sMdvj6CB1pGnlRlKov+BIfqLy+d4Tkqobp3pEXWDMSenSuvos
lEISwXG9NfPvcVWwXkR0okyTh4zBbvtPxLFOs3x5/twDiWe/W3MZA7J9QwOd9Pqu
sJzQGWeBxtUJm/CCoU+40G8rxFm3ldRN+jK34uhQtQgKAkT+3vorZ/PqHlNMNVAF
IxmHhJwJKPBXlY09qJ7LqR5SVj3cC8hOC4pPG8HRtiuSU652DjFbpbeOJXCJ2oBg
usM1wXNoMexyWEunovcf4IXSsMGdcNfC14+hCDR7SUtqCoGkBajx8Ma1jRzVmo7u
12WGW8vJFfBP3R3tVQI2CTCHJ2Ue+R0LfRECNTKXU18XmiQQnEpmKTgbTFG50jGR
fURVGBS0DjPeYa4g1iD536SSsJqaB21mTi27otu1t5RFa4UkVpkqTnYwoTSg9F67
mdJx2rf7LinKiXw1LlJ2LaIVDCl5tvSGA2yigHTTcGjHdSdNMztZ/dTVsGC4TCF+
U5c0ZnrI7GDy6qVociAsFROCSYzD5G8ZslU4G1ZSUB7OAe1LxTDx+hxm3cxxy93c
sKLo6gkGz2aUQaohCSL1GaH1cc43KTXc6/zoL3kQyK9UoOGSeYGZYkS8DKh9Lrdk
k4nhTd2vorfJfTw6Ugtl/b/igLJupZoKzur+jkx7slXMbr4Q3aaxLpkAR5rjVEem
xxPuFCyEwp11Cnisq/TGo2wtR+2oRi3yLF8DldIrClVZA41S3n2YmW1S7h8BudDH
GUrds1QYXVWdKzqhGDUaH9tDYcvIZ+/J1UNjQxGJGR33xaYoyBllp7mc+SKjdb50
24Fji+7D55dBSk0OGYk4ovBWAJ7reJWufznewRfPuJZQ0wPwwzkZn/B/PXEbaPZx
2/WCy7DhoW8pXvvzn8ySbBZ44omp+D6QjhCI0AhfUX+0ajguzbqyddPWeYEEarkS
8xTJMq6VmCrLEQt2E1AMDYonKWWuHGukFm0+NEMFrSkQoxx52pUDT5F5FpgEqM8r
R29qrB52pRxEiO4i82OkzVgLcWgyP93vKAnWZRfIG/HOeV3PtVziqLl2YYzD5Fji
ClPf2daRHIpmocXDtHks/c30DmuQsjPcklh9hMyXCK5rypfs7xzmPDMX+A96bzH8
ItvJTBEKaeloWhSdXgjlruM74saI+pP5xC9XVB082PZj1+Z50evYMBiGJ1qriFgu
Dd1DjWdqR7P0FNtB9ypGzdrR2pI+Ae/d9rxsyVKfcVf9GVJtpK8Jx6JQzj3gQMxl
Jm+M8/SrIxM33/PD3L2nrmFui1bCY0IgydokyWVq47HbTTCHUWVTqApjzKV30vya
TPqRleRVPAUElBDoQCl7GTvuF3j/fNmhHw0bS+mTt67fXVSQ4gkTvO2YFK2mMPas
9OLKvAf3NF3hfj6hzrVU7E3E1ptzOVCY3osoQTM9s3SE6slCyOWwBkJBe+WDs6xs
sxjmHTbdnGqV71XzeO8elWGv1M8Q7xHmVGYh/qWB3kiro1UAghle0VJsnkFViEES
YVoOxbBMYjHVg9IyEF1FOPbybX6biV/scqslvE9pV5e02lNI0prTKHARAcCp1yFq
LkCiV/tC+wvGfGT3wcl0PbuuQpa/nnd3mpNv6S3wzsK91iDygdRVfO3AOgSgREpG
6aUym0nvBECuIqMRyYnWeXgU0r2DBfVxkqIlQDucF9wwXw8iSdH46uhlSsxZgZWt
uXlyK2/G+KDWphIMZCPzFf+NrRtkuHMoxOC//Y2vX2xV4gf3b3Ze0LzPra1Wxxqm
YdvRebWV6Px0NkAAoTHpDDOk1NQAj/2MGiocQEquO3rUe0PJPr2OcEYByYixnJPZ
0RXuZTdIDrrPt5wGoBFPFIhlO+I6Y5du8bBKo41qeERzURcskVQmWNDhymt3CaAD
DhhGCccdn9/wSLVIapEMmsRZCGAjnIrjY+NVWfXg3gx4YsfksA8Tye5G6xpVMwfx
xXhJeN7JwTtG/Uuy+T70FG91HFDXpxdN37TqzogQrwWByj1I6Nvi5uba1njygHcD
r23drw8cZlRj7qBjj0z5ZGuInQIrJqmSW4M3koeX5BegcLDFs54cFgfjHKOaehab
gN4zaZc4v1v8zYNgNSK6PrxDmoG96mAxgTxP2NF3RiyV0ydlN3HkhPSTk5Kk4aZY
5AT0B1LbPJT2qytOKm57zDEdNGGxr8R9EwJEA8goZlDtpSMDcpzAAfO84ItF+SFC
mxI/qWsuKg2j3qPU8KyASyWzX0AcLkBhCa3Vcxrrf0wzs3w6p+3rreniB25lchYc
lDNOsJ5oJ6bnlWLKn/KJ+df1YiE9eZAEgx7VUwc2ZQNzLvXUU0n7x+PshPPfMrcz
nzGgCaPQ7TSM0l1yEJStfeGxvjGA8M5TvzQ3WeSVL8tyFkdWpCMcGnj8G68D88RM
0xJ6ch8Kwp6YCRfRvy06zvse1DRuT66Wc7fekPbAEsLhs3uIZ3hMsllW+FDP8VHk
Fk7wkGvmoqOjdGef72b0HySBIckMrPqLKO+dcd/zb77zi+pA9NxKIR2NnyEcs+c+
hkM6TwtVGnmLcIlFXrgfwVn8fZ450dJJ5cmeVqR70iQA40qlbyM8SDkRkwhyBeFU
E+8Ezg/SWSO9fKhK9lIPucOAK30fUzSHqxWekCHRQfDUsn/CVo6w4ww8VlVKzpsy
cb58vzDGWrshoObYM2rij+CPM40CmbQySf80G0zYye7RNqjhlswdyW/x2baa+h28
LgZM1PjHPUDru5RV9ViL6XmytxLIh0j7u4revIvnSC/4HMAzDISwTYt/SnZ58hFN
JWGQHKIcUui2MskQYLyFuGnot05BQS1ZjciiecaqePLh2o1IspeVJEAtyOLbJfJR
N3YcODS00avNuCy3Z3i7+n5P8CZYxIQPhWUmB/QdciBv9wgofGAc1EGjQTMqzbMH
LoZU1TbhpfuYs4Z1H4U4bPTdEuJrO6C1pfWfBdqFpluWxPDEUeH5a8Y0FMcVKvah
L674UQMBUBxSCzSLFaDbYVNiKHCl8IotONP2AECo/jocEX/t6//1+3ctc2PBDhTb
3saKUoUMz3MYhXjzLUouCws9nnzJ0uBVl07imQG7uYtR7TfQiaoeIhC1yxrLrnsM
nHpE8p0XkXtE0yx0W0Au15dlU4bBmjgtzp/HBIMPK+V/ltFR3d4uQS4TV7mqIdZY
j238Nh3UsR1hQefXaTxcCgzEgHOqOkdw+Gabqs5Osd/bcl7R8L5Je9AKhA3Eerjt
4VmNTAy/RdiTMBQugJ/knPxAsBRMmxMQrP5jHpwf0XD3HjgD00rdNm6rzwDIlO1n
7j3DufBcXI0qDN0Y9cpe3OlOmPcGqhYZt9DaSEKO/5GJNi9M2xquyjsN2p63XaxU
bQ9J1rahgjdS5/MYLt6AHS0ge1e4fxinFdkMHGDfBA3td1/qaYZKWmK54od14tI4
928FAEYL/q5SndR4EkcdG8ufiTnSRhTBM0UjZhqG2peGilrvf8AewSoPNFwYo4na
1HRIH/j+C4aQeZ6/1HSw36ex8ElvzMhyRV1B2YKBOP/ZLHsA2odCyK0PzNtjA/ye
CyEB263tj3cn581vm2nQPY4ertY0OHHCRjhCoSaNJCwPKDRGYURXopliUu/eMued
XodjEIiKuKEJ823CjbKpBdHzW45VozDiN4KNS3qbbg7G4SJypV/c/fex/LYMDNh7
zpWdjduKZrkuLe3cGjcVqh7eImhIC4MZ/NmYM626J1f5Iens3vrUmn/tmPvU0ckB
URkmShlBvDy5TogVwrGrmvGpol59Cy6HniMtMbIYf6fNj7f0hoMTwtBoQvs18faM
TyPFPunhyQ/GBP/2KSc10iGUAjJo94k0n/4vqn7d2fLv1BPZ1jo7qXBBCKUGkJu5
/F8GBncktGjA3qj+2ZfJELn1mROQNpzB3qG+wvJJoPRsV30asGaOni8mtOPGEHS+
YgRSJCxz9drjU/cg0n1goMnqdrBKNIk/1y8aAewagBTk7P35h4LNbL9yJB1uOB+N
M4OtTHshWtMpilsVyUO1gF3n0LxsdZd8KBDszniZR8lmCAt8UW7rIaNsjV9NH8Sy
jhLjyiCh534kz90g+75hkyNY4XgdNoXO2bh305/yjpiRhuRaKRZWYGPm9Q7eEHer
9I3I65R5Dln1zuevETLe6GfIqWwHeDFEvJvLRUjU1alkPTbCdq1cN/Tyo4sFmsLf
l6D8VjmuRGOsfH4ky9CRUvlPMt0NRqGkrrNgA24qNvAzKwMgho3eN2D+Tj7e8SA4
ppG+J/wyxQrv2BEC5Psw+E6QaGwDeBQj+AKTdnbNb2eb3QHu2jqnlkRqHnSyrzM6
bPKlvG3iU0dfr/yFWVGgz+pmq+Ua2ojw7kPmoTfxeZJc+CgTVfcnMdOalhbM1Ovn
yWJntOIdykHxImmC9m3hXn17754Iy7P/xJuFCfcQOuqeLx1C8+VRg1GVNE/Yf48S
MO2r/dMZ9W7q8yxRM8eTG6KUwqK8Rz/tNsip//sKMBXSVNjmao+rvCK6F4z4mDOk
aG7WvSwXnO++7koIyyvy/PAEjl9OPNAv6M42TDl9JB1Zm+7goBYahQlxWk+/b5uR
iARogAm5z5iXk+W8eeiByxrQetsGqYbFWnObpIQbWGOvkTO1qoyWQZ6sZiEqbXNl
fW5D+jXCOsx/G/7ASyKghtFPINEVR42HKOBuUBFvOeEMlpike2S+oMnQrqUQCiYG
Y8hs4ZBL7E9saU+8ZS38nGe56U2t+2TYB/NZrmXouzY7t5kxO+00aSTGclGctQzh
wM2sYPO2XEt1UF1vUL4sE0hC91+mKIitfjVHnmQHuhrwNXLUuLvJzehEDHtxTrLj
nq7GZLeAhm2p13d/aFAGwcKs6BoPPS0wDMxkp3bCkFC4GtCaFk9SXWHoUIOPhZsa
+/Tc2yEBozrKQA0pncJBsWIXWpYftjtel4E0FqMnAYwYqGLvQiQfPgNlkxTp7dvR
Y8WwOmC+IzgQx63GGWP4qE3zumruscJvxV6UeBRfiO66Eo8kD0uXmUsxAn+wQWLF
pfQqpP/bRgnhpVMyQNvAQahSiCTHXA+xI/90Y1di/+rqC2QCPpih5jFG/BjbEg3e
WYLvEfQAogwIg2Sm9FBCpQ9QOJZOqTpW7Fjazd5Z1l4MYZquQ532xoFHsR8wrbSE
tV9ThCaNOyUj9lBxYaOb1/KGy8yL82Qr9AaldgGOhjsqAyVBQXwTcmNWNZURv1nF
TXVcgTL83qz5y/KzYPxaVfuXsM6iUC1uybJHAJS1RcCvWYJwidaqVJxZJ+iZtc5s
ws5RveCEzmbH3J38Fyn4ZDI1PHaVllkUWVyPkrzyMR6AqYmfaWrei5dc/ZgPhHNY
MuG8W4e2EKzal5UpTe8W2Go3B8aZa1JtxJcg5KsZqe4nGHxchhaZK0qpRrcjuky/
rdhDEfuOS5WQv0Myqa3/5rw4VuS6vo+DyzP+DrKnkCX7GzGwd3Ptqp9tb8f0e8yu
5FJ01c2Hf4HyP298yb0gXbfkLkcqIhny+0WlyWlmLgLaXN2KRsyzD1R3RwbxNOMk
Kxp88o85h4ZL8l8R4KWbxmEM1OLTI4C2z8AoiWXlSqYU6GS1nj7rgwxiIbLEsSdf
yD6I5umDKsyfnUJ8UArVa2EtCLIZ6Oe/V6+75oo+6yc5snT2ZwsQQTFaGJ/8FxD2
hrA9INS/ZeC06kgog364fM4dIps64uBl1e0DgqvU/+7xiHTnm/H/ElazuiOxWrOt
R88ytXHYY2PNMDG7xHFEYoQ2ib6xpy6QpHT4tEY696y2bDM4ERYJfkKj+UoQ5Jzu
JOoEBmoGLLeyaXTB9EUY3U/ln4Z+rZvfW8YXgWpxXpdQicvY8RFlmi2Z6mhynupT
qaieSlHTicTZsi5iaee1yevDTBueSK1jb9kymgpsZW9aYWjdJ/lhnn0w/KHUxwZA
395mPsjd4K7BU2U5FKLkTLzeXMbn9iTl51IfrW4a06ByadvhJeLKh36pTTa2fGJe
qqrzr7c3BukAr8NKZdAuwYWAZytTeR30QfGIdA7tSeR7jdRJz+4HaHnnzCgIRsy2
G/0psOAcXEJVLBcE0Nimx8i0zG7+6JTpWJNi63xPIrYHW2Uaz4SidrYUH6Ng/kiW
CKlE5s7jzYllWJJxx3OjaBQrDkpk7W6LTGLA2zd5Mot/TWWNZSUUaCdi6+dnRwc+
wLcU3KlLIBo/ZQlhu3c6dURI4kOkmul53qJff4rGlRFzoJ+DNeqGAc5JONDcT5ep
aKAu4qhTd5197n51Gn+6FENzrjVvCliL5/Jy9OuMUYZudmPF7uMP4JUjIWqODN10
WjTplDbbh9IXty70xA2nzBq01Rake5kghZe74KCBdZpVs4jCwXrLj/gWjgtXuQKP
jG/utsDk9EEkxWpcE1bIXesHEvljsF41WAPjzF22uVh4+TyLy/h2+7RwhlN1UPyZ
SCQS6CSOLh21FkLq2aFez7hUQehkLXhJFYjYZYMisoYJGsQm67ew5u6HsVhUzdht
UlHAZnNIumyEG10bcidzp6T7tebTBs6VEA5MKf+yJesrayyjATEPfiRHrFU9R8Vl
bAygo6SY+2bwIRMClrxeBWrQ5WHn5V7cBSrb7O5dRsigGczY6kkTFrYIsw9jftOO
j5cX9KcD1ECLizJto1bSuNHaZz1UVJ5suYtbC2M0AkNtu0rrsC9xcyThKX0eTQgY
TSqrkWj1zMCbFqBLIeYDFuFbkjt1XtF4h3KC28wobebpqzgKynQE+ZDpLBGIXZGv
xRgUe4XV1LNIc7hBO6Fk1uET4jvQZTil71nFWOTa5nGEBwFsP2UHpDgSX+bxOOU6
nKyooiwWRPkuDlpEBQJ1NRcBiwCyYJ+eX7Xl9X3GfB4s44AxMG9BmUmNkMAuQcF4
6VeFK9I/PRA4tPL1/JzB4ZZj/Feb51ZVSlUWLH+P8ufl7Z196tCMxlFH0vp1HR6m
Ya/etwkfYdyHuJq2WQXOz4mfO3x/azb1eoj0ouD/LqLhR757EbiBv2qKihEahtL0
/j2ji+lacR02pE0c6aKL/+MRp4lusU33qtLnX1zFfXlOpemoajvYtJeFRi4JkRxb
fCuCHv/oF61WODD5fZdeZdpLa+qbqHPblgumc5PQh7XOPLelGHt/q/WzLpDpFMkm
ySFBbSVldBpPAVGywLNxUV33J7BZoh9/3CKXRYBQGmMSU08gj9NA1QeqNmfyFdJ8
tti5aNoa6rrPtODt9aChtagDMPE4Gaebteo6Uy3JbvPqACuhm36mFzOZyuQlheDW
Eti3ZV7tb4gvGPfjfBJet0vE8BpE1lThOQd9JW7VzTFSfycbmXSy23KxQPZ3hjQj
GA14ubJcPXweWgirsAs/glySd6a4r5CcYHMlZ87pg+u5i0clDcyNt8/Gw0HPSEfh
lMhhwaYekOOfI+xgHJHXhWF+B07yvJI6uyn90/YgCvEs7a0kxZJUq2Jf9Dh6vuvy
FdMgalM3MGJfp/sIS2pTBorVGWlg0GF1w4qNVeaVvo/g/+au5atZI37b0YEDtObu
YLrxP/a4jl3CPC2ScBk9V2JJc9Whc6LBnRbXmYuXIa8cBzEjAEMCOuCMONcEadUK
yU7Ch7aPqXdNi0W4GBqcFXVDkSRhjySY1Nzwm0SDwfog3PP7DFBl4Xv2kjUmWlvZ
QYOOkerTNR8SfOGcRuz22UjKpPlFj5dVFzVeLWyv35RzTx9uqsoo+k+8E2eqdnQJ
bEnGpPcfFRfKinqM7azIE20kGo2SNDGaCJeGjUOqo3Dh+3G8Y1koQwoqNnLCdzYC
34s2pBS/fXXc4OP3TOfT8KokTivydLU8cenJnASzcj0xru6b6sjciWrz4FXlg92y
tqN8MPEOBg1mP0xqV5SE+ngJepAUUCq3GxbEZc8M5UTrXEAvIfaYyHBZ/9lUUBiS
rj8dXZcyIZvgROLNXjpMb5Rry/qH2xoL5jKL3COrp9WiUZf8fSZrhFoY6jXBmi1n
bkq+JhC/Kd+rBkP4NL/NH12gNd/YbfMyvaVdKmZVAte/FCaMrI3gZWOysrC7f3uz
hUnxr33GQVqm10WxynN5jsCe3JcvBKl2mYpt2SapF8jwSi/Fta/m41df7TaNKg6Z
W5QryOyFTltsafrF7Lw1/Az6kLb2HgUCx3hIWbbGAAb3g/V/Ne8Ue/eyNk9oOj8C
qJOICJsh0TOu0hlJG8rCw8RnnKnoXe/LkXZkrdcYoZvTJ0YVM0f/aEU6LWdNLlsI
QZvsca7NYJOov0J+7FS8AMc2LX8A3AUlQOjUeZk1b1dPY901akaifAgEeUgLJa3l
pnlcY6rnEpfxwdZ50bDDs6vbYoVOJqckwxR1IjWPWTepTvzEEr57eSoiXFNYx518
/u9VfaEnUUzrBr3ko9eEUQ2c+8mvVrGofCGdHtAp25UlFNCnIRfdu/gU1q2R0XlW
Aaa5ZnYWrT5M/d/U6/gJpfyKZKWisAywYJCtu2Pq0jeVzb1CnkDjWm2wEdJzj7IE
SVc9jUz1IXDPPgnvPZz2uTyAN0DugQEvaOt0pguisOm8AtdJPJ4bSgZcqE4jd91W
sgfsIH54UJOuYjf9td6DESwdUcT7raqz1jSn+KSx2ziRHBeCKqr3sL+XSDKNHrjJ
HpJJ9WYeyXd0u4ig3CqxGA7a1ThNKh1KEaEIVy24a7WWFpiNX6u13KOQEaUSljuz
cZUohCXN97gHaG3yxNpcc43+KMwm10HupSB5zRVBXMWk4q1AMiNddxeNGF19NOxu
YkRGUae+OiNlFCvnfnkqOkYAvDycbyDSR61FTIA0kPSDa3nEs0YV48Y8RMaHJjVS
fjfXomVZpmUTD5dEND0qaiz1MaJxsS4TQFZQphUWkGem/4go4/ZHWV1/WMp0QaSM
OzmlH13WwKxhfGDFDkxDpW4fpf9lfd7uX4WZvKqSfYBD0RZ0JQCewBqlCBnPPA84
T9I+P/eAMngctDnc/6NT0JR2huEpBps5BZVt/PzYu4hrMt68uX0Gc/UwpaNLdzp8
FEN2OyERUJwNSrw2Ly+Qv9dEAbVe/7HVuHN+c6jnZ2lPQcZOzFn/HLZqwIXyYvL9
3vXhjI6tVQSTpG+j//Iqk7vwSrlbEICtD6AG2/YYiax2ILQjlEMKvD8LfObLJHG/
xp+AyBOtORMK1XtOUvBdjW/BQveg3G84O56GueFXrZIrcn8CVjgbyBonieGlBPtH
Gzd6Uq3nBGostXIMZnQLI+evBLHN4IgyNYA7llE3dKnMuw4zXIT3gw7NyFLzDIPs
D1YyZtlQGTf45hDmxSkkKltOe64GoUgwH/fuF+EzQsdatOotQTs/ZgySKfTPPnyH
gcdskNe2DczUIeXZX5ELFUbItAjou6UmvYHyVtqW8EWxbaOnZ06ro5cKmQ69O9Gy
Fz31JSbMOSigDSyBKBIixiIOe5scHzG2iQ+kyYVakynD85rw1MPCdM5C1++wQ5XM
uQKS5LI460skXErTV2JIgA96f0GUQzQzKIaf29iwemh1ZTOwaqNHypdNvsJyUcHj
RsAK6aP8t/b/yAQXtCUUYRYtIoTEQhMlNZOp2m8Y/T+WA/BTzNp2WMJZmJvX2HFd
mn2/A6pLr9pY+6uTK5vW1ad2G3KsnhKbLoWTQzV3U+ZY18YHw+KNQT1x1pCacQrX
6W7t2dGbQqd2XoclR0U17A3KplSPeVSgqb4XVTsQTmMlTPwJ6BAOEDB9nErP8QtB
VpHvYoRx1iRw9MJyNtLEHiQYxmnt9cRoFJeiN93hHRpneitexCQVgStqkMBWjgvj
Y4YmwvR1PjZfPMhRdH1lv3MbcLEXBWOFjG/HHvWm3Zj56mI6G3nvNlUkQVllCBOy
dWEA1PZnen9Z0ziAWnuohximm114ZFXBwc8YSvuXvlDPshPP4D5ji5Bvk3CFs/wI
Fdl3JG9pCwrNmHSM2wZlY82gTXJu0vJKFUB4YVsaCY/AHaTWFjanCroTB4MXgQRj
hpua/BowKBlY6nMezY2yUtJnHCCNOscm9d2NfWbPJbkxtgFdXYZSA/okqzxIeDgQ
4rDqmuhJZ7F6e7Fc6bMfOtb78x7bHEfetNwU4dIG5rLG5KfAPL1Ns5lTWfMjmb4W
oJAOUTZq9VPcoWuA83Y2vulAKDLixCZF0GurAgTJXPihsjtlIoIDnFvEIoxG1Inp
PLenSciJh7srlbCJZ2XkSWg0uY8yHXtdJQ/7/SiNOamvRlCV0Gkv8cQsoezSfdFD
fRdieKcZ4WRxm9uxGRq3whVDRsGGqZG85SsSsPH6hhXBl2srtiK/sqSg1Es3t+Ty
TWVNVa0UOhYMW8qpA6ex33fxvMGaqlUyPR9RvDJnzogc65IlhynL7CfxvwukqAr/
CQmDyjCQOHT8tkNqn5ZO5W6r1V/H6fdtI47Du6+RstpLYsl9+G7UjNYG4h2a5AdT
jxZWOWzbLpfhUNqN97NLX1KGd2gXbURx2z7MAThrkmngUYwtH1IE/nGIjsOyF+fr
hmKfDfDakk62+Gz2GThyLL4icugq32wZ+YVZH4DTSp+EQJDZE2UUiZBrhrPQXM7/
niG3mutLLWFypvZYC7SA3i6Z9O3Bzkmn+wQVVTvh9zPNsqp3xwen/IfppnkliwT2
KNFliW8as732esI6QAIoNC7/Iys1E7YULOcRBDA4SPvsOTN3ZeDvtDfVfoG3YE1W
vO/0QE7+WwYHGHQ/D5XlOFiXkCmpnOww53y3dFOGLgoMeuB8Q6KFt1/yiHx1QZaM
LPlnISCbY2dKeszURj9O0W++r2aDnIEI0AqsIhlKRponCA9TxksoDglDjE7zr4kH
hat9xVpiIc6nLnTSJS/DgCr/ZHGb3+hQ/7Fmg7K1r9nR5r5gZWqgJXCRJjUjXE3T
OaDxzUnJdEqvPg79Hr9EZQLlT1p9JfD6skyqZyvb1+zhUcmshJfUHNoWxfGKIyFQ
0Fxdlq/3gvsWG6kcUNeAVNwMIsUk29QyCVOnOaKJ2RElWQv7OxzJJxC8HNL8FWzb
isLjoo8EjmWMYjFrmpjrR4wZBRf8wdb9lHSu7hiSYI3450OEqQ/zNVVAIQbOrHR3
T/STNDLFM5JZuuPKq1Jvv/9gMdwO5syMBvqunjz6P5UbMOEhmGlzBTOtPVrvi2i0
wnRLFGf/FHTsqKKkQ5YEGX5HQ+0auEP+A+CsY98ct95ORHMYo6mKwq7Q8nuRS7ct
EVijPtrJ61wqh4y9kbcoovu/TjUR5MZmHWmNRzMz3EGjmTKxt6BZLyQLEUys6vBR
PU+yWPUre0cnyzkgdguJBr65lNY3UGqSktU4j36fZKznEmNaZHolg5pQyBHjDbUH
FNOFOA4eQwepAC6Xtdgh+ZYyJssGY/VwQSKxT6yr+fcd6z1DonYw4JKr0ZFC4mix
3HIb/qORpWYcLO9OX8uDWlOuPi5eOFl3KKlyg5VMy9begcCbcMoaGmbg2dxKJa5S
u221v5KNS24+ZvHrXwmkoA01mrkS/PLQ22/cNUv124Hj1CmwD5hqZAA/PbWl/9Rl
KwMPdAITo/eoCnjpxBYSPCTqhfc52xk8w+GHOgG9gduCz/YKRHmwZrBu55G83cgO
keiN7c5bI4BRJwmYXLqT9k/wJSNlHYGTMY7KC3aPR1dH0b0iS+32jOXWWXnyBAKy
GbI+El9vjVEKLSix4jGSb8bklNcKCx/wPkgpQjs0pRx4VB/8ET/Aa47+G5/h2OBu
Jq/sJ2hKCOXcVkAiYRrhV/vt1qwuF4A+BUBopK76FeF1Zy6mkYiCgEv1+0Xr0jt1
ji4ANhKNtTLdqKl62heYUUMcY3qXlxkgH9JWPeU7EfnTyAO/OGnvGLFatvBRn2Xl
zvmmwyaeB0BNwmDSR4LdiInMUPbTQud7RaSPmxBFAGp0Df5RWOnUDJeOo0J4aW/L
wkq2nf3u5vA7MgWbi5wXA3kLnt2sCZmluiBKKUnxmQr1zy47W7e4m1MOXgirCaLH
rnCnZad3uVX1JV03n21Gjy+G6EIxkknWtrK7ML+/5KlTrV9/zh/UQheSJTiGFnsu
Fsecnvgnm1z5xD3Q/7q6DD2AvGBhBiKguZV8chIo4xSIXAMnoretRS9rdJ7U2FOP
JVB5ru5y/Ayw3X7E5hUdvVChJiHZk9O8GsYmVcAetVPQ9n+I25ppqWu/seWjG/de
GPuRgs6RTjimw9nnX8X+Jq6PZ0C91tRKBrQoMDmguqI6TAcDkHtJwEINA1xen5bC
2/i1iuj63IK40ftwkMvW9ApxQFPTzSIYv+6ReruPTUPXH+SpCmFi2igvBpZE/u+i
Jdq/k9X1ZXPAFZka5FX+EgM1UHL+Od2QvDBKbSrs4ribMEUehH41hU/Abg4jQ8jw
VfX+/vthnX5BUqOzsmE/MzVbK89EVmC7ajfIIH9VJ9d3BOkOIE6N9hiWXj+Q0kNV
vu70c8/E981jPkriQVm5RU8UTwVcPDUV3wOLlWEcTka0HAuuXHf9JmlenfaB9tet
V9UryRTTN8lf4B5e6LWfZEl0BEg/cpvnRLgmXkS8p+SELm70PaX+6WAmH6XQfRch
qOLwrUL7FbDFJ8ECEyZPffTyAw5VbcbN5omg8+UZHtmXAb/4OX2ciXl84xKE1xIO
vTwSXIjKoKaxrjRQn2ExyHKKW9EtrCjYwhWA43dV/ZFTl3jEhb130Ij3sMMGnAAW
oApNwPwxS4sNrs2+ZdpqSvt80VCE1LWcCMgNGpwWa5WS+Ao/WzqocAvc64rHzX2g
RUrqnDM+6g1p6NuG1agLw0BItSkOuZaOPOUN+J5/BqL/st4xmDkkCoZlnI1eXSNV
ALW2QVaz61vpGqzaKaTGkyvQAM8THrb5fAEExDXaDysh+N1NgqX5z0I9b/G4/hh/
oUVk4KyDKgDBQ7fTmqg1JY1eBR+ndw9MLXWLDRPIUEOJzZQYqMZ70faMddsVZFH9
fbQaDfSuv306qHcU5yf9dyUusTTxZAivsRGXnZyhe+Ylqmz1N+nU9wDrVVimzErx
iLOihg9zZzHy0pN92T+B+Ix0SHZFN3u+UAS437lxQoji5bIqTqZO3TKhjnqr9/hf
HiCZDje4FpKFgwVN9DOrT1Eb8Oyp0iVSWAmq5t4TEsdFYpWry4yaUAEoezemrbPq
ekygN7H5KkerEgdECuBM2F6Vre5XBO20dZVA2UpO/Nr3DsZXcSH24SRi+QMYSzhr
k4kxgRGop9HOR3yDBpLzUFeUqsycfseqmstu/phE+sDbi18yawB+wZhIEmDwzxN4
gIJlVFPwCAdzvUB7Vwb+j7TCoDALNdtEv2vwnUa9dwsAktXGYPIZ5cee26XiwGfT
Kp+E16NjBe8QRl/jbttqXRY9D1idmgUsWjdFY5y93ZyCRqFGaMenv8BvMHDndx0Z
mfN3O/m7YGVzj7aTfqIOL/CmxtjtZ1luOgm3i9aAcS+mtuUjnUkzVZjmrQ2NTc1H
QJrAOU1wdFwMHQVIZ73tmsB6A1boTlz0DpU5Q5ZlD4L110a2MMb/VFSyJD/JKcvT
pKf/MiUQyiMerw25XkZ6JoK4TB53RGMXAAaC2iEcsiTFShCKvZlUlfQPI81rtZon
J+PvspvBD7kDG50YMc4LdzuLRrwQrM1LtUuCGjAIySgF2HlkVzKMjNmSYRE6nsbX
vVAghwOOjZAdMmzXhBKI0cLD4yc2tun+WChwuEpl1xHtzlnY/LkyKSHMZQwl3Tzr
EV8rvwJQ3HLZljELtYh2dmDFLXqfDCGwbPmYDwzY/fLHSq4KvbRxC7FtiXcTpvlA
yOW7zTksbcn3RGKW0KDq0vATmq4qyR9ASsCTAauklpHFkYlUQZn/aboW6Ymw4xOD
rfyN5RKoQl2zVyMzSm2SoGCea9Ky2SDl911f3PSW0U50H8iwVcy0ATCHjiFy7XWb
5IThxYMh9Wf45Oe+NQ2vbrFN6H135ysHRXotBDDxhQ8z6HdxwOsjrrjIOFCWuZU0
GzHcKCRztFyvPc0y2MZT/HFArSaZN6EEZgE+k8IsHIzKiHR6NFcv1z3jx2FLZCVd
hZypZ3j7y5H/StcM/RATG6TjgJo4eHL4QlVMKJ9zc2+YpdzGs2F6qe/jky/KxX2V
ywMDIELxcMafPFt3HUVYh5aw0Y+INnR66sWA5jLVEnnaVV7tJDRZEF6TxBYl2n1A
VYOjmyUIA8SJK+avCskFr//sfEnTqjGLrcIMHRIbU2pN5cG0bKit02f38RquC33/
1O9JcJOSk1TtCEyvOH4qAww0VVpLWhJaF0ksJ0sBYrAhKmBL8bNfV8W8v3oukbGV
alcJlQjjpGj5bOv6IMKVGTC22/4GCLQLh4kVHEGtWFBy05xGJrAVnIaKA0WbYaXT
ldvWjylD6OxKxlw/HSWHRIR5kvBHv827mjpwiHg2aZWWCa3p09vms65xe46Q01jL
wpKR1PYXNlP2pozoNZShfDN+wG7PIZnOdLePm9pb6peOh63SEyAeaTML0h0d8BaU
xVot8/sWKgt9qxkB2RTmCz4i82J8ikFIrcuWfQoTPbQV2rZNrUd5lIHuXzXLFOwU
cJt5D6kqwEToWw53LiaNlLvRNTKsNhBMau3rVp4TqQ65Wbeeau3h0jn7OM7SMTy4
dyA0CGUMrktqiu3tkQe0OBz2MSpcAKngyihh7IAFnu5Mrh74DIc5A77GM9JZcAhX
DWLl+bNEQM+j/4ZnZkUCcmwmYcSlMMXQetY0jvmGuCCa54Era7yny5UpZpR2Onps
IBZ1W0D4e4ndMMvOnsnHMx8wfn9WXVjSaHyJI+74Posor3BhV7eihb/C6jJU1Xpj
UuSioag5ciJ2cxAhLL402gZi7/eJDqpvJQ3Ht5eJoOCcE8J5GTMDqLehVTW2pvQP
GRP5Y6wBvVum9QrX/a7Lu1unp0hDdpGCvuAs1MdBCR0+IGoDhxGEEbMP6pIglipt
coBrvhMbq/50YEazRSt7dg4837UYPWKMC7kQKpRpl5twX5XLavASSIsIUh99AOcn
vqixAivD6/KVxRoqZ9jp+xBaQCYbS5lt3PVaUl/KP6xkEzMK9P9osX8eIQgnI0Ok
zpa6T5JEh00K33JE3dQb+9YuZts/Zq+Us7RY/oWcwCl5jiVh5dpazG11X/6oKMDX
2grQXrDzJ1fMJWwSlkZGjpjyUonZvb+sK6Cgyo4/jlskCSBl6VIBdhIkpHG9UvIQ
3z/vhHHHwCzdhc8GsxLyakHpMEelU/aI4l5ID+T68TmTybebGd8xb1RHAo1mkufd
U5IFonsqeZxTt4aakJSETLg2YczenbfRcBnq7ZnDE5Z5bJNcfM3/j1Y2Dk6SqpKb
c1wRpZzWE26C+d6EZ09iWxntIGjh8J/KWrRhGpRDG1rl532Hghh2lv7svNibmA8g
Gcj5/Vajeu3phgoNrGhppBjW/KUkxT26E/eYT22uBbtDOPFMUHUXYZkTqEegdpVA
0Px8wib7O4pBuZlHyrMaJ4xl0tqQutA/LZMpizY89nST1pa9QcJ1+/PWOUqlZkaS
dPTDIDUzBHqJD3fuDndl5F4lLeJYwTnk5ChzEh7HM8MovcJgLYcK4AKlNnBVnOfb
FN0qDbcS2ruM2LHkIUViK7saV2sZhP21pis19O8lPenRRvOxKZWt2YPF4SyS6+P/
FTJnTk9ew1BdSjEsGr7Kyk/kr1OGmE3t50ztbxPq2OgG1DAvFqCJL6DKmjhq4AG8
S5fIgX9MGUqLKyT49/HV2fj884WK+Lyhv7Iqw26Y0gi+ZYHcQ0H354Yi77c28JBb
WzSna2raoAK0x572PNbXOcPSATtbfruKo3vQ+jnQ7DqEMgovs2TazBdGT0ct3FMM
Z6OFI11+9noGoPy/ERCQsN5OQ/f2f+iVD6wI4jm12QNO5gKcWtx4gtbmXV9D3Qm/
UZTubOrx52qrm8QX9xNtoAuw9dATLbySb2ScPPp4GLXoFSiSr2pzt7jpYVreDy5P
6YQvmyNCvOwPfftzK7pnnCRVY210jQ3n7AeQrSO+/aVhW8Tnfy+aOE2FetpkZ2gH
TyUkghpPoEHkGXpIPx1qJ/Zw87Zd7HxiWQTdFEQxH4LXrbvsv+9L8Q5jxlYUHtQI
ZDkyOJNIEyevlGWpnEMxjsnNtyR8tAZuMWbJGRfLE04IRpXKOqd3pTgkgeltYaYc
yEW2lBXiPmAqind67UcGnU1e82B/fbKFqbfttNcm31ZZtebgQkaTac2VLqA6f165
xNAkpFT0nlz+x49G82G03bOpF/ws6SFAAMDCq1fQ4VzWaR8kc2oeG/0YYRvvr8Da
OycpisEEw2WAEO0OCFkRnDM6Aas5IJpPKd4QPJDdh8KFPSEmbyow5TlR18GwDwdL
9v4ReJOFZ7BAHjc4Rw1CGvLEZS8iPJ/8YBm0qNQi76obDrOzXEKKaIMBZ2wGfj4z
NzwpuuISUroemUT3XQMo9V7Xzx+VcZCLGrzxH9smsDIDhpU/MUQG8rCWKSBIsFeI
F3Iggj9F6iKfavxal2EGfi0SrPNJRMDpMEScMVRkDknLLqM0xvgndtI5WQanHVN+
QUyZGlqcmMhf8FTwx2Q0UZkqp+PB55QcIiDHrNXP4q/xpynXWuo6i7hTPPCVW0EG
McWeh54gzQPh/5zG76wAwOq8u3YzGN/40jkhG0Ce224RauzpBhVBpBWN/I2D8+6C
edk4UlAWwO96bTQhxuiDzCUEHZCwrgb2InVa45rAWI7UXfzCkYHhDcH2Gs8QW6cH
ib0zwhzKuh14idd3KCQZybBFKcb++kqHdpgKzolQCu29dxyCbiv7LCQoev72opzI
s+D+cxEaFHqTAiFvWUs1qHTEiDyJOufCgTPoWYFqi+mIEVnNTIyyn988aMBxq7Q3
39fhVfaSG9XS+EBgJ068uiBITq3slBvlfzWgYQjyBUMN9yive5ndJT3M80o8BYMk
Lfikix57vtBDMHZxmvrao99jyiObXX18MWHipn+Htj2EiiKnLUqQwnFOyrbqVktK
MMja8WQlRWHLc7Y+/46ab7rSbHdr23FjklxfqtbD5ecwsCD29KeO928J7ZD1CH4d
eHdDZCXzbx1bVqXdb8BjjizLNdN30fvFz7CTQHzmJluySc6up1c6aBNi2TtbXdBD
eyzS2gI+ZMyUkgE0NR+DwBPliQT2w+YGk2N6P1mT8VPf3fOXP0AR1Az1Q7pt/3de
rO0wXGTmJrBNXOw/qg5YavK3fJjYWHsRZIxPdICUM+PGNgJ3Jmm6uqMaR79qaG1G
4bz24YMw6oG2ukC+nOdRS6NYF7X4UjX/hhnWGhN3GtH60YQZTMAS49RE7BhEP/kQ
4bJOvfYypGLGxhAeZf7n78wmFeB+fZacrcKDkyqVTTrLEKGknML49YWIv8VFtuEv
ZGpudZXh5zIYPSjw6vUHdQIj6NSzuLNsaxp5ozDSxdNb1VpeWd/ymUk3DNQ7O5fM
oKpHOSOTWzvoAUU9SckGzRNasT5lP9uaU95Yqv0yc5UT9kUbwzjMx6ZK/yBu3Hz0
PF9kw9cysg+SRF0OiMzLM6glyJFAzOvTwwlBiILBS/RrlKRuA8lYDObaSaraDbEd
QahEf8L7GcBP9k6WeCcGk8GsSCYqWQGFRrZjTDugSX4G9mwILPta/zM9NiulRgT5
XfOI6Y25rpBY3Fn1X7aPe+NwVUsOuIieH0W1jH0gK1OFXvptq20UGveRum+Tl4aP
E4yZKSy0BOzSQYruXhLWteirGW/lMbWFe3O08gl0svfS8oeENhA1NAJZhu8lWbIK
XpLqpZ3WDNf2A+hOi9/VVgN1IMUZxKf3rGxSx/ISJXNNI0lwATaJHG8LaqgQejbZ
iZ4KONUs7rIdGh5wB75+Mhij/7vWcpjcd4X414VVwSBTso3QVb9Z75/8R0rUOy6c
onLvLxlnLtI0QCLnEi4Dx+hHiILMkzTCqeOgmQPw2ur+/Uz6ahIiM7QAxkpiOROl
TGl/vwn3MKQmT/A1JINOgL5WpNN69ZYXjLELFtkX5XPfNG9Y3E1wSDctSBncEhW1
0ijqLo1+Rp52DiKvoC96ARue/4JwBpX6niATKDYnimxN6QWMsnB8VcUbNt5x1RO+
mLw+AyXQg7+KxUGy6LjOsawVAsgTYZSFCHimqPzSfxnefNfqRLsP+sKC1q4Sstme
blHEh50N5JSk+m7RkbN8UDtHvGPDXQg1LWKo2eX7LIEqgcyBdIRKE6DkBcGg6Ct5
ETP/Wbp14+nrzsvCaVIctrCsocgQtjjlJVNDgUBO7g7/s6lFQwJFX6eCideZhs5G
TtVnl53/fjO4nOqAZL0SPyxV2YE3wlOii7ybGXTEzg60D/d+RHmKbefHhiNUAvtl
yyyVLptZuuwIIentKXimd0gLMSgZL6MQ9ZXoDRp1+/pohxHvAa6cUKYt4/s24qro
QvB2a8xdHvllSJy+NMEOtqPqb6CZDCSjRCiQh3JMcocdIN6eiUnA1pESp0jJKDcQ
VOuDnkUkxi39nQBb0kdJbBzVVYQOJwQZ4wa2u5uUmu3c9GfHKgn++f2vrutj6Z1/
XJmpBktboA0ENTladHGeYMOHOwErkOY2eAVLi8UMc/A/6JJ0XGIEerpcbYWQsWLm
obIi6gEOd2gBkE8Mthr8K5gpoGbSEIUAyxUzjOH9vD9XANz/2iWB0oBhHfhxk5T5
0FkYvmkuayK09Sg3a1bvgMBSDJoVBtPtw0EeC9ucSAygXmvhdFau3z1Eya4I70ZT
+VTAeVq7/FFLm4EHyunEFRt94vaDtW+UIjoMx0CitxUnW7LfV8/UhtsV4mqCRjsz
nDbbLW2/hl1sUtf9YeXGKyRRGMEPl7trc5tENqoeEW9hr3dyFdqvLwV2bVWcSr2G
mR+gwj8+coZCVYb+GRLesfVVe42i4j3XVq30wCFaQZh6lYs5q6yo/6Z8KpzqWMb7
MmC0t25Fy6nRt5nl6RgNTBsrkpp1drJIZjark3rmc1reD+2igiaC4ItA2cWwG4BT
2jRft3vdUB7DBVoZOf3LPX89CXLSd7LYfNxRaPH7Ek8jtREHOxtBwbLCbY+4V2Xq
f0GofkSGda3o9OSujJdewggP1fu+5eC++DZGfiyP0vu2UHhx8nPmfj2RqYeId+l9
9HPlxUNsAk+Tm6zNJA4qlldXeklxOtQp8D4btgsR96H9ibur3ifiCEnqtw2zv7a5
74o/5ublQ3c0cPoIzziFuxHTCgigkr31zlJ12sFochKH01M8JjKW0YbZqy/j81c+
aXHT6mzuxEi8/2P14hgd1yi04S/VRUd+HlVkEFc+iREq56YNtIeEfpL7YYMGTo0k
K8WEXjE+wuWDD8IOjV/gVozxTZ5yABj66PsYv0yQ8nu8C7x2TtDeOWjSLmqbOTYf
fhlDrDV2UxWRM2MVHl8QKoBj096B5qTTMhABK7xz6miWL/AnJjg4CAE7QWibai3Q
T/e5QD4M4kxKWNWq988P5/GF1lMfUqcMO46WgZV6vtaUdytDNjr7JczN65RZ66ef
sfbxOCHmDGkShPerzz3/G6dWxkZARI9axeUPuBKnLjpXj16FytYy+adO5nQbOjvO
UIfwl/YxmCsM5a5NNAzMhmxQvsRt+fKtLweYqXz5ranfquM7tDJ8G2TGBNysElHL
fuB1M/n4VEijWBG6mAF7TOFb3O+j2P27KclginKDCcgwU3vAoMiS7s8o/69c9+SD
kdPKB7jPvsPcLpWN56aBrNIwkt3skkvCcWBiKoxmgco8otCb/oJaroEPamiNDiTF
4wy71Xbjwo6C4uRrW1NLB214ki5RpSUCHEDgFO+xU44IHouYdGJvHtvROAnNHtJn
eAyePWo9ytBXrit5NN5jxDbc9lr05mhWgSyCBk92pD6Li5hf27mcWWArRLXRTqpo
IqqRyiNu/cWNGXdYp8ymxA55v9stU2jexwQiFClNb90hdLnnPJjS3IJ2UmP5pH7m
WeSP94ag4Z7+xfmF+LvSr94CQGBX508CKhcriomr9hPzlV8XKDY90NRbUKpKiy7c
D+aipL5QAlNLy4Gv2b5O2EfdDRDV1BfTpWhoTrJ/OA73P0SSvqA9X7u2O1Ps7N5A
sa/jIgx0CNOS0fA/TKdnCjqGDtzOsu3soGBx9Du2DrK500gkNf7bAKa1+tYDsuge
6MK1Eqt1PfVdr6XW1603PgSVFivfjyLZR4V/BdUipYt8GN7x96ji0caECax+QiS2
joz6viKo9JlmBTY8BWy670NZ+qlgLjGI9kmDAnuPYeRQ8rMvWuwTsFkEiQPJTt51
+YOea6qfbniDjnd0Ag52o9wz50pUPgRw6pQJJJ1uTxPwVz8wBM/xrxtDJ4ewzM9j
oo9qxc7KtVX2y854D0xO5GCtTrWC78rt/BF6M9sJtByBVY17263HWWj+marNHaul
ycpwLRz+fEda8D9NU9sR2BFBskwhZ+wRVcmekaHx94dwRjcQCUiaJPXm9nKXo4V+
XM6zItnJuxHAlT2jkzQBbPZJ1e1hZh1qXztQwycuWRo/3TR8alrBoIF5qHER4tIR
o+1smvliweCEihdAvquzHSabVTk7n4lXhR19P2A1MOy78Zw6TGNewMa9wVg9thAm
OzNfK0dJGKd1h6GKNABLcVRfmyU73CKjA0CBfTVTfvIdt7pQi0o2+gJxvP6xuClP
SdzEPvzVuZQxu/r5nzhESKdgOUBJXXJWbBl5bmp74wP2mNmve5G5Hj72tScFfYF2
01NXPkEnWEvN1/r1dI8kdqBmyvG3v0Mbn3QD9onr9HDXTUOk4m63CAyJzmMWXt7+
sziYx7VOPHO7po2NetSHtyXpLd22MlXtcWANk3knKnEctz2QZO+HjSoU2D66/1M5
my1Vcl8dg9gdeHBGsqdDTGItWc7SLvmgCA5MCl13/5WL63lZzTR1bk7N9lY98OjI
FQGME3Jfa1x7BEP7epMmf1eXSftEn22BkXLNfyEAksMO1O3ELyLqQ8mesu9ADNNJ
yNKuDDNKWk2UgD4ZgxIxhXpaDx1Rm5l2rttyYTRiIC6D24MHmm3OaOUFzi0VSfkF
QY0BWqqyCz5XuncBIUsWVHX/7F7wJEaImzatrKCULs0vGPnrdYNG/J/CwMmXgEC6
VP2RM5WM0cCH8RTeo5ZwJezxUNRwtW8sxMGuqctVprxNdq/1FiN5vGNc4uFHNol+
rI+utLUiWYh6NQ5IB1JOBEr8z6FH7n+G9aE0KhDBoL/aJ+6cG9BEAGxdQld8IaAM
zSWnylrZbES1vkJVb/vgwdTJcWoC/0t5tP7/kY8t9Cf1+w5BN0BOFl23Fd8TPp2J
8WUnSYhne3NhygkJV3Xf8fDS0UaLNSuSe/DbUE+iprWrsTF31ms2Lwt1kUD+3SNr
i3o7bo7Fzi1T1qO0C5lQpYA6KMJZnPxswh8ZZcioswdtywfq8sCV8a0Z+Bxue+Fy
pav3Vy0bnB0qQaVWuj+e1qC1cysRejxxDxeXOma5hSCvZVLZrPZGD29W1FzYh6qe
Kcpa5yIFgXVwQp/CTuFcB+I6dHPtvPrSrOq27rM3JMNxvXXNOuUK8NMu7IVRAWEo
Uurhpn0qCkfqieGtBJpby5PIw7ELNBYl1iNhIIQkayv+OasdRL9rejxe68AaTiHc
1+uPR0px7rfcvZLp4dyNl81qbZoB48C9qpq63Mr1iruMNkzQ5cYF7a7pDHmNA38Y
vC0CyaOjmBDFf1dQnqsut0LK1GvtzQogjBubsmB/FZyiQgnr31HUH6aAJM2EA/mC
rPzEDOTUxF603oogMeONEb3QUCgpV2moLURAsqjI0A6GQmM9Pij+V08t0/3Wwugy
KEwRgjsdBfVG+IW0UWKXzY7i2BGQarqgR3RkokPAjbeYZohTLPPRNdCo95yjt0C+
3BsbvWqIcKpDJzBuwmwuAfemxgdzREBoqJiyUJl/1laYwqtux7MII/rSu0vvqcKl
cQDr4CuvVERRSs7IrQx8S96kjOY+nDNs4Vu6Z6d8B5fudWWOAHP52pGvwXd5rxZM
jVRM85Bo1ZXUIPU92YIWN8519Kk+pU+vrC047bKXN+qUye6rTMDet+qR8+5aMIjq
aseqOsyeqXbFyQIwFuYgXpubrOBVdGuI2P8BMBtoMAjDHO+gqUmVJBUmmuYJs07E
q8QmVKjy0f3qEssTLuQMmmM/smZO19YLueZeJJVmrMm5sZ+QDNaWZtOp5II7lXWH
Fmm8wqjwpxGCobtx11StPc/nxApKStdDOADTsvbhoqwQYVksfgAjkX4AR5QPrO87
TXgwzZRohqNIgjm5LFam1Q7jZcN23wlwQ7qi4mGzQv/xt2ej3XNmdhKlR5f8h/5n
nfHqetogeaxvj8HWJ+MPpNlh6E4uXdd0TNXsNDSmyf83AqTDi/BuD/EZylj8Ei2T
LBwuCnUC5Z4zTLen1mDXm4uJRxrnSfqMxMJd2uOVPWKw7UiJuPa4XB3pqU+sPedQ
q+Jzka0PYFyxY0Fjd9+Cyjs96/o1bRQLDxfyveXxjec7NtuDj+xO620wKlwabFEK
mUwuMEnLH++znpbwZJZGHxSiBuLB1tuJBbHR99jo0F0E4vLbDPP0PjEbUduBt/ZJ
1fs45j3yOJIvBZuNY6kVBJTcW8ha4uKaEtiUIfj053QZKzFA268KIAqscoZDutQ3
enWiDZTbX5r8TnkVgGLvWPOJPZ+rSnsjuITVi4cvgbto02rL6pJyQNC/DoPTKPMv
PjRNOhIBB4gT/bjML8amrcgueSG9Huhp3AsSGEuZUO2L6EVgaYCcO2XSwa1Nl+sj
MyIvWZAB4OaZWFIcJixgdi/Oj2iBeejSQizdvQiPZTb1o4PTR6cmUWh9p8rvvZ75
Cm2ZHex9wGLm/cCRdWq5o/sZwn7QAGCx6zfU6EJeF99IUlhsjcexPPEpeRT43Mfq
cjCvClruIPuMnKqAXLzNfZe1oQdDgzE/9YxY+QrMVpTq3wQklmYLLKw5IcZnkQl/
m+h7lrQ58ZI5qLGfd4O6fuNC2brr87Ghhi0ggyWNFSV7LIzNXPr0duLKfHerZF2b
rbLbi45WViAJ+p4J0DTAgTeyTicpVXi6iijYujww3eNFvzaAiSLGuYVMaJk9zI+0
sq79MCVX9QyTqBKj9kGNYyiZgjtLUTLzACysRvZlvCRFutH3cL0RRwr4vfi3Jrln
rTuLnKFMqqi9hCffjiOb/1JSF5P/X/KrkBbG0pvRGgsM9jlu2bWjMnDnbbSd8G7x
z15O8qrW9QDq9jolfVlKdATZ3oUWBGwv/qa/R3JMA1R/syBvpXYqLOeEHzzbBLTs
d0SntbXL35zr1+5ZFv49oy6UN+Jb2HtGgvykZi6QGjwcKQmdt5xM+of6YsVaIS+b
YlTmv34NByn49Y6t17EwmcWv4aIpf9JDbePiQ7xW8LCabykN9+6nVRX3vFzUDBto
2VemFEdcNJ7+bEMnTEq2mVSZaYyk/Cfhp3nDBKF02XHvAiBVOlrZh2sx6tCFTz9l
wNcKcnyiqhK+NuvPIS6P8367FvPxrVznY6xL5AXnEn2NjHkiNoZ3S14OaSGmY1Ce
pn+3WJa6O2Azip8VEo6LP/Hc9EpshUeuKGZhS+ye/aDAM2sPjtmzsODxPihGvHbx
7G16iYNcysHkCrUkKayuDVlFN3KNwjGL4K3ibNMGff3eMj1piG/BiW+uSwXEbNh9
vVUniMtiNCJxN/E0NOS8xw3mIs/SwG1g0jSyffVRHvz5Zhc/o+1wBLTeDo1WQIBu
ZdUTIomVFvOPmJKazGZ8+OqZ0XRG/tAVZPofRJ82pNVccrdtmimeOWVkZHc9R8Lk
oFwfCtLZ0vXiXMD/JZUGcCrWO9rEswXwXN47BHwtr33xm0phlGXKLZ++rWMnG+XR
iZ3K7BoSsy2SORMRIx/Cy/iL8M/RmMSCnRQdM3rp6nhLwkyvwU4LJSZoxYf/cCQt
7HFXcWX+GXKGp6apA0yRCpZGy3Fm1LAyAtuvFPr0pme4nIVxn3F95/AAfMixWPVa
TcNfUGFwezt8BNTtapIu31Kw63bQbfbQTsaRx29mgOTLKPZrqBI0r6CKaH71WN9B
qNqZFAQ0ot459ordcnZBZZkT7MotGHnN3hcBrBtuH4zl4aaZJlmprGVE6Lkp2aIe
/x+WvZiay9vJJo3JY+NaXH3coT8SY+lB9O736Mlz5jnFoIkEpTdPpeRqjH0zE89Q
waDA9zNVXlJ/c6wkqB+fKs7uRcLynV0jHXpi3acXgE3lU/sXvuSQn302dxf3hw6v
H3I2MekgdmXR4ajZPdDKn9nnVf26M0qt3hbOio+tdemVgRL/qLKX5KRgleyOdp0F
cobnLoppYP4XcvsUYuATPGCDf1KnYmRSnPriw5H7DdMVf0rn8623TB8AWbZr8Za2
uY7Oil/VHSZVasLaVrkWzx6JajKZlOmP+5uPGPgCMfmCAww+z6gPSO42wPgATlyi
3h/Zz6m0K/vL0CPudoaNrO/ob7wBr7EZXeg7teic1MbV+Etq2CfGgtlJjY7MvP3s
ixkdS0tMSU86II9+gLuDqmO8+OY8M5fSY9L4wwb8LnA1XE5EzSCxKvNDc8+4jkNS
PTRiofRV2oHBiYNOuHjitB6dHSa9Fch5gxd3eUkfjqlsKmJgcKe2MllMmMJz0DBc
FhZYJ1VuXIVSNlq3m0U8gR9s6h3+ANbyXE7U4I/65YRylzuSY4L4V38/+UVHKLDQ
O8AkYIqXCxIc7W8cKBreX4uynHKjW5z696IIwNe7xq29IbMP951XdknoaGzBejvn
y3SsrlgqqRQpDNlRU0uPTOPjHXlHhQDEoJCOkYP27i7KsfdiKVHuUpGmQ1gEAAQN
cs1lNsZFphPn77/zCe7skFuhLLGpPcwoelqRIpl/zqxx5yud7EB3oYDQo0sBSpWg
L35vxRuCoAHWQ1lz2roTnFvWf6VRchT9RMTR+TboRUTB+8o+fouyeoSKJ2Z4Nem+
0LI2I3DV3hOvPvCzUr+pVdNjIcwdjb3vA6VS+TngGe2H7OdC2YywKZFV4vieaJLA
DuBnCNSkbwexzvWpm5anyMWTRkDSgtcm/rQfWGoFow5SkqS4+j3VO1CzhQFlHVv+
9xyXu9wHTJyBON7N+oLnNCcyVe33OKGYX7LF1WtE+e8ahdhEDDUuZdceGCaAC5xa
xYQfyelpZX5lQ5jzY+PTWqpXAMsabLwpYjqlVaa8yWOyXlBDW73rqFTosV1Fi5WC
JBC9Qxh9icPwSFKcDAYpyOoj6aTrAjqSkWqKavAE+Oig8LfjLJ/34UU64AApmjmq
k6dtekjN7sWAgUVgLzU4KwcWKxabyqi3JL9vHvGe1uCj9k9A6AzV5NjbQB3J5oXE
3km/Zeg747Ps3V6kKjDoYppecq2GSlhNxXBNJBsh9Xoi4NHukOYMu/nBug8aniN4
8GYknFALU2zzdVQe/QiQCSlsgqZ1UqDYS8e5NYUNFH/JY7ri1A9m9hL8ZTWbnjdC
lAONLZK+vXv+XKwFHHW0tUr20VyqkO7/ICkiXrceGxQESA/fMlaZFR3k7hbNwvZl
xSfaJTn7TiHzzSB1ZiZR3bIN0nAXwaYYmZij2l+cZ2Amd2pdDYQI9q11/EmYPozj
vjG9zZdc/phEmUXNZmLVeJbG608nOlTVsbdtKlxn5cC65dUP05YpRY4csE5oDnd6
oDeZ3lgIztDSLrnGQXTYhgLEDjdbMfXgddB/HPFlaYYCGgcrKsCcf2VUiEEFSQFc
MPlbg7nwKKLR2KG+sVupPCCBRHFk3wjG5JPUwMuk8+I2bZTGdhVz8Af2eJzGZUAz
kGB1sv9N2EyfhpeE2LHvB3hlz+lbMvA0Oj2eL1q1XL0UUAq+UU4Q8jiRakAGOuQ6
PJ6bbQFNiqmMmkGWwj25GZhC0p/dUM74PJSyEgnDESLjOUNpi1QtpyKiYHKftnbc
FU+4watT9M6FkbPGDMSRsJYkJfXzeFuRt//WvPdRADacqd97Gz0pULw4YgpCdNqa
l4unbvKrhV2K7N7xj2POqBN2p+DGbqN2L4wRTbFpRErIHxwcD45IYJgA4StaEHzX
B/ZMWoM6+juudX2Tc1LEev2+UcufGmGG/ZLAXM+xG3nzidfYh9yX2p9Oq1YeErXy
1mAlJw8evxiUXlH+9QaKf7++AsBWsXbrg4JiWZYrcQhRcUgOHNH3hj9NatBrKLOX
dF20B2xZNm2ljOqmNFNnEKGq54cL6D4RzAvkcoBHPD0yWaqYlday//lfg4SElI26
1K+yG5DMGZhFpSjPrmUIfdSj/MW6Lq4ic9kJ4SOIs6dd9+iYEU5AfVsDHa8m6z6v
iBcC+hTN/K+kENCc2jhlv/BC3c0bLKxK/tf9AXXihCOKGG16IBMTmB6Gv9klTwEJ
VYkOP7wu9j7cXYxrK2IOIhBwscMfQcBJzBnOA+fh0sb6RbN5ID7ynDRYAATgMnh/
FflP4AH951ZO6mEu7vyKpMSHPE1UX8YRiOlFf2vTKE5tJ7uuq/FVurT7UCUBCRbg
rh5i/lsQe8OOLWdzERCQhwRBfZ9ZAtz7ra2DijEtTz8uC2cq6YxP+05HlhrUbmR1
7/FDJY7PIB9fgcEPnBM+fNuWwm47Pbl/iAMGN7vPKwk0/YE3NSAxNJ1bK9h4jeyu
TxY+KOBS0IvJFxaC6S+5ySumJ6LNQXhbuSRvK4fgFHTiUmh3PIfkiur1jI+GBvuR
RnNXXFNRBm+KyFUMMY9shXyBrG74oDSgNDZIXvcbHmrpBXZqHd/sAM/2lqnXNSuo
ukFB2vTkLI9pernXMeUnoh1mfyUGUrrti3Pwu7izZHEjLgvGUnQn/0uhtQ2rtxiD
r6OH5ymk1ijpvLn+VyqutMBJkDzfGHsrFyekwtiIfy8yR+cyUDS2GRL6bdMgx1kp
UPoK1M+mIOgd/LcI6fIsCYDRW09QeBRXJG5NgiIBYf1QUbpaSE5xerSkwM1iBN73
mbrOhhE4dUwHdsxn0p7otkLlXKT4XCJJpkNMz/0Q0k/bvZjOOnFe+JB8W0Qf1Ixb
zTOj4sg5b0vgCTyGsazA0kaQ63PaCoUsRe1AyaG0dx0NPLp5Bv2gNFusWkVbrV6l
21AXA5DkUDh/vGgcNxjLDLRMh0JmIh6V4Jl1/EnH8hQD7ObBUTnYNYs+77+7UExl
brQLa2akfDM+ElY3BFR+smce7D0i6tbetbB32TdbKIuh1SZtXFE8iB7Pf17SG8rr
tBaOb2ETLtyyUiB3hfRFy3j3OGKbUWb/84Y5dwqbu/yL438Pqe5L4uq40PVPXN8L
h068O3LhpK+vW/PsIshKG1j2J8jK+HvWQHiMDV+UFOGSj8JTzyUUcK994QmK/AvO
aKl/3zC0DARd+KEaukCOqEVwAHFRvxAE9r1Ynpps7PcsEhs8a0EJvcNunXepJUnX
zQPysynDiPvjBbAWdEjwRta0SufIOpmGUpAQRmISOQfe+CdzHOLUvE3BD7CU67r7
1PVwCtAJ0CL84zjXK/Kp84sFrIYkJFL6zKgJ3S5mUfgn1urZ1mhlE7iVqw4MvVG7
dN68ei+E+1QJFmxin8cdFduNTRdOZnk+l7vvD47HTyLNVFo6VtgCd/u86YGOzUO/
th/toPtrD8iLozCXnj01lZBYY5sSLlqismjN/ZEtioE/SLZa35i1StOO7d6+I1hs
vfcs58hla2cwAfdCcNPC2XYvH+JxzKjc00o17cdHun837OkQaLlmZDS5pwim2FnT
JOG1uXFPCh/fhH/3SxmqkLRipmIjEcWf/oy0NiZlVB/S15IaLzj1eheWb5YjfhgI
AEsz6nQjOIqa52eSgTgviTiHV029tUc073B7mD8Qoi+YCSt5ir9seFjoxVJlvOl0
lQNPd+esdfdGzExj4JnsdwJOLp3V7lZpFx/tj1aNFzxf76z/GJzoeLMWkDfssD/k
fVSvak7rEr/yVTEMtpBVcMIWPIx+ckpDIJq26svLKVgsu2Y8pqEE2mu4Mqr7aMEt
g/NkYFOr1Mhy0RqDp1dhl61jBwisSkHt0AXsmXXcI6KuSfHgJeDvXZBMd6iF0WLX
2kSYKTvHQ9uowJclF51b1in74sdjzeqNF/ecSN/MdVcRXLmbdt7CtQXyebxpqNDg
W3aprDyhEty5qP7pTUcOW2knHR5xlogyLFCXS6jNGU6nAZ4ev8nUmofjKQ6Vakom
wLVBpOUlwUU7EZxldADleiNBv4XaN+XEmQS7xJs3/CzPqvThNntDzqD3HhuKwmyL
efq+CJs4g2aqe8b6HHQMV0AgR1AJc1XGIqN1MiCBytZjniszlh9ltnWMOqQXlScI
Lw+HI5hfkqH+KtFehtxXMn+avkkNBqMw75Z2Br93al8zAVG57hP8LDJk6plEYi/g
rC0AEC5zV5z02lGsaW2ahowYvqMpmti+GWzXMYBJD7sCnBHolB3q4jdzYsCrNkUk
oRFk5GDQmb5z6sAC9iy/192Gmqetbe0IsjqbyVvr4I+/gE7aXOnKDo22RF39nLeE
SXrmJAOgQJ53xpw0ed0oRcankqYkC3DOlILguEDQ/ujHxUVyXcn8EINysnKxhQcD
Tf8OX/2MST3lkkSnDwdGn792wt5H9T3gHXs0057MVLfNHIn6fJ8EsuLHP2AA8+hd
OrbBJZAzQ4mhYvcEdb7N/R10Ud0S4gtJduPlx5PX04FRoLErhFnbpJTqV7UcmZM7
4dLNUoC0e7piSOUZ0lcFDCTRZ7Q+f3Sn3g7WvvXdStwlAQxaOYwOF8thqLr3o5dd
jU8RXzUIa6+Xu4+UUlibIU91pqXn/BZQtTCZTxQQfcCNMH/GhOuG8RapX69IIj7x
lR5vYQ7MOq3MC0cE0kVjCaRrF3MIIb3797zkrGSXBp8tlTpvfm92ATXcjqimVuOZ
0ZI7IRwb8wkJDUAQqoVcTDIPlU89RerQKKN2AW1sjbHEXX1NZ19p23tb+be4wpPw
HJW2xIG0+HwvvPXDKMzlhgo9et6PIExFZK8ueLgEGcsiOwYQuRrhttzRliAtDwo2
OQB7KucGdTwLKIlxAKmk16c/olHPXTZtN+ERvRPtGmzMQLP4uusz3Adixo6o1V3M
9exYnq4hkwnBrkjmBlzrco1uxBiI3cq4isFIYsBtdDV2dh80m4VxnRMUGGdGkA3x
RA+1ZC7/y+t/1GqE43WJ21fJLOpy25XqdJuFDPlj2WrWaU2Inmn3bcbCyiUMlQiu
7/84eCxJHai/E/WxvohLFDmUpsepyT8vymAs0LIV0Ku3Fz+HyiMp8k8eCXusGMYR
4aaTehgszglqTn2FuaEcHmFr5PEXiGClbaivf4pqz5ITrEKX4qmJZrhyVQBKajNY
6ebyM76x4fuSKMfGYF2qS24k0DIFSrFi52bSILQ7MlKRJ8/ziPJUKKaKXEwk39SR
SeCIWXE0222ofDEM+WsbmzoDOJFKiZqyWTI+a62t+JJyDVyfsWKF+hFGdgvpqyyK
FBKOXiL4Tbg1BIDuaniRJwDiOofoBmM9BN7ORwRwPx4FK07+mMv7DWNatB+6uc1u
+lkl8BqT8aZMrX6YR10ozVabggvFINe9ZkLizttAkuVEk4Dz58AH9k4umAIJ2huU
ZcNM5pim9P1ZhOFYdk1sVphQwHSnOPwWKCYAV9BFEi/hBHCONyLyTasgExV2Mxc1
DJ4Ixu4GW4quw1fuHDjQIontaNr/XTB1AxDo7pg5YwWsjtWDgXFJPC+mG6O9x8Bv
hW90GnqJXgHnk3u+J3XRifdcrZT9m5DXQZgPdhED22sbI4/Pg04m2J3L6FQrNsYG
TH45BhZRizoP0AHVq1JqDL8Th6aUsu2pUMVDleRP7VeHGq7vLCSxpQED2VErLPLP
IgWFUEjZYBumTYbbdoMGCL41xoMvHZUr9B5kXPwFHRg0t8TIJTvxAuaBzHhAm1j9
iKaGvU3Iw0zrW8pgY9gKqhCabxGO9x1SU7c4HhiyYB43MF6Ir4tmuhFoYGcyDjHD
haBHayo4IXdEMEbSwb/wF+rqJRjfZ5KASyLx8fRSjyzdWnalBYopIChaa9iIO9BH
L9WPS6T7vveL6qUZ7aF17pFH9VGU4raxvxK5AQkVsCr5eyR82UmUrfW82EQYNbv9
NURRPtJhNBJ/u/gZmQMbZsKIfDDQPhfXg+06xUKVKPDv1Jj9I7TOxBPpzB47WZ5s
BcGNThwJS7MvqO3cX5MotQakuXPS99P2FRYSXWlqEBg3Yepy1UPNzL8goKIN4dMd
4APq1HK0o3OyXeaqc+JbmexxnKpdfcEr2WuYecp5ibWSFcpFKZds4lQcHzjZMe+/
ZFEnrkvx49siwKzTfVNYfgaGysDEE1wOy+DezHICW8PDtAqDP5clBFDIpkejf1ev
pbp7C1hFokiGzMOCA4fo8BWBVANCmJqw+NfqCnC8O1swK1wh3ViB50dZ4Q1sP95B
XrCDyEAB0jsw1sJ8+AjVlS4tUCn1od0yoeqTtaajmkL3ApJ9JrICiNVkfYmvH6Lm
mxXctzTTf/hlAQmNZaJSHJCik78IPg8lLcWJvTUFQMNsxzip/yWPZKJeIVie80nQ
eNyOBT1BgJgfGBX42t7gyguptZqAnlD+BYh5lGa+8TsEooOZAA0ZCFYEXb+6ec2m
ie5guQdnpUc28jyRlunrrcepVS4vq1Vnj22OEyV3pSQH1llXRTpiJDNZgOuUQOXc
e4WVX4a+u9Ry2lO06vQPEyQZ0wCPPkReX8xa6j9+QACvqz+/Un6/N/Qv4WZC+6Wq
I2LbRQa7Pb8QMsFNhWatC4VzCJJszu8YIXAc21CfYfjGC0Jf57Z4DkCZ3N1YEBnS
PawXkdgaykT1n/P8inWkQm/51Y6kHvPJyLOWCCI+0VkCZLIpXxGFTTU4uCD6AeOV
3YOedjm0Uxc/LSw52lklMRXQf4/abNymVlUzAwnB7MiBAGKd5HswN4J87kbtq00C
UjXKy12vGnWKzHHpvdl8Tc555o8PZCNmzAvM30a9GrhndZoZ1F0VOwc5yPoMTQrj
Zs6MXGRyRLfhKTmf9acLJHOWy0DpRlfe+Adk5UfX7sLlGrw4zMQwKUUKP9TOvQxS
kz8Cn+eyE+cJapSV/n4PEo2X3F+2GzM1pAIkvme68VrbQjZ+U6nVLKogKj7niNPE
F1+cCOHOatUNG7U1TQYDWuD8YZNSEvPQR369KIq4+k9XwHFqlV6SdxIto7dkHmQF
m55dTLlHTGo17JLJlZYHkUpcoRxtJ6OFk1Qv3Fx5CdQW+Jql1sEN1gk9E9rTN9kl
TcaT7huRb+A+iUyQnYDpX7SIfzuw31Kg8ztMlaIZniIuUOdYIJy50I4aQ/As0dBd
AqZzvwAtdGoMYb9pDlsv5C0P4qTHzokkRYxOVWmQAuDiNiCu7+h4zuyXGmdu//49
r3UvjMHk4SddH/6L3zpyUt45hWC4g70eYog1US7aiddhoSBPvpaV00OiSRiy/EJQ
KwDMLzA5L7JQ+Qag4ZOg22xO1j8ReeDBTpekfJtcT40NKPST8/rkm4pO8izIU1x9
FnpBzf9gSDO26gs/Sb4GzyjJDY6EWSjGTcoEnbgC1b4JVU2V2fGqcFrhj4Yagr0a
vby6kEIXR3+m5gz3/kEwSM5YFwRH6327n65OrFjbxE3pmfjjbeD7Hza45yKaBLVB
a2EFNRwdbTkztFzSZ3Lr0KMt1DazhfJcaMz/d2FDLY+r9xFvdmcF49L4oM8YACp8
uauBmS/l46K8BU6vzWzP2k1+jEPR57maSaP4pgZChBx/c2NfiozUfZtKHwmeLalf
m62RgZCoihJxiAh7FSQmmbWdulKRxUb8FQK7pecq3Xl6IodgJsYCe/ZXnwVGL3iv
70pwxgZuA1P/lNr1atl7t+SYZ3JdNcif9th35mU5k/JpACFBqSPdL/DUC9IYgE8e
Z2yjC9zCp1OwsY+OcZxaOmrerfMPPu/3QpU+hUz+QpoMx9v7r04jmmk0AsIGL2nk
ttlK+R0ukQV9FLPH+MJSkKLuqFGOxvLXTVL33SxePy9w01irHMPXoomU6I1XO0wI
n5uAMosxwUsamA3QzxsRLkDFCFX7Dp+RwNuecCMcSULD/AYMCGkMpdhZCok5TUnt
wtj7i0E1BHoMUxOslw24IxjZZqyO4+CzgmlgKb/PsC54BF+5ra5/FFCzGIDaqDHs
DFKDNaqLnDpIYTMEYmdbrhSSlPvyp/ox+RnQz4a3ErdYYfTKkjUhb1HEqxzA6F78
yxh+6PauuksPw75zE4Cwyb2YEfKgwuUesvXTlTZfbY1srRoybGOxMtWvBM8pHHfd
DM58TupnyZxjNNCnyRuerSPM7sbCBHfkbjU4qX9iGzdgzmWgFgpCpb1sVuO66nfz
wqSMewFGX/88yVo2dAeH/jxG+Uyq+xfbjZQTQueWg8jE0pugyQHciMeAvWS2J8HM
tgpsPraqty2Qy+4vWJSHDclzHwLb64pCrpkD6b7zJ1Fdurs+tK9vYk2UJ/fTRPWx
CMGGfUP/KicLXs/qQP8CAnG+Ce84/IiBzSOWPD/uqE8uMnfW5u4QX6o4rI7CrwvG
gO6/go6UMm3c6j9UL/q4VXz6oKfSRQvAbm14e7HxdlnB25HgLDssKF/0OlFFCXDT
KkVtQeBV1ylxOzoMQsXgkx9w3FJ0O1IgOYIIo9sBB2lB/rpAsv3sAeSRH64Z9shP
SC4OaatAI8hTurysoby1I4WO1jj7JxcyGlX/ur4r3LhNvhjHBExCbTiOnkuW//j5
3HCnIKdH9K1stfa7VgbvemYltvYBSFpQyrf6oGq4Qg2UHPdRbzifBFgWi6mFJ9OL
ZfjyqlLuTdO8f9QLBmxBKtuZ+oDDXuCSFO7ar7boyWkvz7hhXTBpww7Ifx9sK21s
yPrtDHvsSjK5cxQTQ08ECbXVq7M4tDbYuxnAGi32J+F4o+1cgt0deiKAgDQQsTQW
Qczf6Wk7nJ3UvsQ7NjvcZKvQL+BttWn43vZD6Rwy4sb0IWXCqo1Ek1kDPNQmy/j7
hOOvZtOGVeFqbgKisJxU1a24Gbxawv8yaqKWWjR99bEnKLvnrOo6pM+1TIaW31sT
jiJuF/acxo+k7FJAmoW9WM4miqcftGC1f1lp55+fXEtS9P/wfIp31e1AcDSk6NUk
h0zCXEy1FG7tzjTDS+8PA2OPVD8V9PHEZeclCAgvrpUmbh1t910Ra71rR1e3Ey2f
HUpzOqCYOo3HS7CZo+RsRkQ95aTnITKOKUZiQCAdNwbJnce7bdRFs6PTmO+tympV
Lxk1F7gT/6EyXK4na2RK9b62tBq3edn9GGsrVKbMT+uiaYxPLnrrjwAnK5aBPKU1
jkP9a7Z/7vgUEPaNES/6ZnQrNkFn7hBWGVLdkNNVuo75MNpYu3SkSOcr6kMqGFQn
u3QH+NWNEFdmbGfd6/bQsxcoRMD0QPKvn/ZBt4lKVValf0JI1jbxhUmeOSjZhWpH
fGKrpRubnlrr80uuDUEYSs45YWNsgvD9LLjip4eBbnjq0B9aA5w0TD5fJYs3jLG6
KAfY5ZpOcllxgcyUxW1xSJXLGbaBmstxedRKC8rAhZfKXI+iU7LTcmoVWKbuOhRV
V7rFNtK1IGS6Nhx+bQvxgFgF1g22TJcE2Rm9O73/yWLEq2QtHE346tmIctrAj3Ri
bmkPwExwsxDIJFypz1bsgA58G2l++Clw5Kon8ZwEjsTgd6uqz0+gssi7VIOlUoc5
dNCzBqbzw0plxfhN15j+35+b27PkIhR/aUkOFPQvGZrzy3YTHZUmiGjkn08QhqYQ
D6c7icJjnRmZUvL4OsT6y6sOf0XF/ZXpJGK96o42IzqwyGGsdCxS/iQ5ExZVxLni
vxJgOjlZcm1AGg8Q8J60ZOxRzJEc3PBypBkQF72nlMqQ3pCnjsvxtNu1Pui+xHND
9C2x8ye3ja/b3xZIUfBTmKUkg6BTcbMeESbqseglM6uKW4jWCbHA3vOI0oF19KaU
etgojmuTOVaVrYWmJSnsyk+EqOH3v+sreT2HaKLC0lFLro2e9SAZ1kDS5c3qcun0
RXYMFOCikLHUNWgyKSJr8gCmDT38vY/PEGJGhKxMrLiz+rHMjukJIwZb3BCTg+Ud
a6YzEnsYQamUcZmRVjbf4gns+vboAQKedF6g6uoItbFDpg/yzhVqhNXXAvF/VIMH
aOc70J1B5p552xBfu06cuxHinWe3ALTN0DU3lP4Ixvwmkc15ZMwyilsdIqahFpg0
9p+2I6E8550HRrXfPgv7AOikZq+VCCAxgUYgCwrB7QyM9xeQxDxwf3BGtrHkUBoB
x6qPwikFV6l3wzToqh3AtN/21iY91P5jICXqTokbZRH4jrSP+jZKojqWFcKrbVH9
X3BaZTx58HDeCR4voTt+VdZ7ZpB7rcjYs0kL5jzUDIuMdgnveMDboQZcC98x3Nld
PPWfI0xiYSo+aatGcb4mELX+n6VQvZxjabYrKKStRK6wNJvhmntbrzjRyvcrJT6c
NyqnFAh32PmRXP+qgnFtKbqc+p3qAjq7B6uhSheCwNishEAELzpRAPFAY+AUFxDn
jMOcJc4hAkjRrWa4BeveHaM15GQWr05OOlQnz7hLLMHKWXSbTs/OiyTFL+sKRbrC
9KoT2EmeumI+z9UP5fPjqICFEiW90ZmMeaYtBlzYA8JLN0f8UFrb7/v6Px/vbZek
2B3f5wqzaPMr0Dc/MekzEWkw/XotveeSDc0KCTGjk+7rka3wPHuVwoKh7mlIU2oQ
EeGQ9AltHwmDUzgwOOKmxj0AQMg8mMjDLZQZkMKMazv4wbb6wrKuU/J1YNn4Z+Z5
GoQD+1dXDrE6QYWZAH95Xc78cqjUFX3NFjbOisjbx9kDld29+MuYTpmgKPR+yCUW
kWVcmDW3Vs2bA9DwsiXkXWyUEZlh0RjVArz2fkD7gdNDgMosubqvljTA0qDydMrv
VxfQgq+7TMKhhkep2ovWkmYgpgNN+faT1NclRe0/bze1/sueyj7LxzQqjPh9iWMo
W3/80hfDwQ51j31J8ZkRBStqArFXlplw70NAxlNBVm5GPuKlfimW0qUUTQeDS1OG
e7mueS7HTxCObnJw/V64LRpniNrYsuPh4BkMwn8a9tj+8J6Eu+atUHyS961TQ5hJ
HxPEgJn8qZJT1XfNuyUXQFf50ZqVw5gRDofL6jNTBeOXL9qK7Ka1C3Uw6VoFiVEY
rtn2Lr8bFxpVqYAfc076E2eiDbaCkcnYplswL6C3qobdCtikSVM9znHl9K2VlwIi
+Y7O7BRPQLAlwmQo4WKwFS4Q762l1ABhWdMpy/Ywa93kV+utv9kFq6Hyoat97my6
kCXBzf1Jb6SdrNqbhhCfMpAFvn9N8V56fjUMkoRZH7hF0y6jDE67CTyzxmPVxxZ6
f9zR2jFiDGbhYwnop7p3JG/3cvXYY5G9hVQvQzELo+RBF3C1JSmLrsqk2GC4TvNl
7uDBZjhohafDqYaPLXLGE/kXAaegHkRCug7vdTqYb/6iJPbCsm4AVjfC6QEB7Rte
Bu+Bnf3Oqkq2KR67kkKHGpaX6DFwt64strg7fh2UTQm6EnhI5R2aCHrIvl6ZFyie
qUgW+r4XJ1Fl9jXUiRMQgj0nNDyMTxkLItqGAKCDlkx6DjL+3det2aNU6Ij+VArG
T3k96KNgwGxRjx5cJqX1RhE1mTUB5vP66RgPdsBPldpGnoo9APeUZqYNfdG1J5qf
xUUQNlcnTMV92+aUmq4drM0XbLG0lAw2Bu6tE21tjJH8FUkckhCQbOivQxRLBEXG
8PEhOfz+46QZ8l+boc9QqYHoA0n6/ns1PIvmqVWphGG0GquXd7iyYzqSUx6nalEg
gmg8N1SzSpMO9eEdNyhFQxhp+VYU25XpBG4sxYep57+Q4Jlh/9z/f3vXYjXPMp3Z
Pej/ILZVP7WWMA/U3I2cRFRMXCnE15K7k4iQBK9bAMuB9kzCty/nQ2Uyze6q3OA9
nGzKdw0qOS8J26z0YA4wKkGJzh+AotYzMD4gFDSbT5hCyrbaZ51hJhZqp0ppl0br
tFpYZgtptPjH3h6RGpl9fiE9h6Ql03mBxEHTq94OHC0mnLKc51bzcSt/tZHUvhbU
22nV6Z8LVGLq49Sutf1YT3fOKinDrhqEJ+JaoAdJrRdZroHVqxFxAToe8wZ93yHG
nd7eb5LoRfFJYU2mPzbZ9Kbbv2EsBjvPysfL3p8pQjzHEDrdouLN0ve2vkqKZqmD
gSuAZSGrIe1z4PBIQ0nKIvq+ssyIke1ZMOkXhY3YC59fMrgGPR1XTSvI3OC34Q4B
bzAs50HoTtjgElaxCdOzqVmnXBD00z3sKGYXAZxRABQWZ63HTlsIo4Zu2sElEEFM
NjCT2VMyrXBt7bBGTzCJinYVlRSRiDGndCvSoUMOHk+L93bnkclhi7SBOGkd3zFy
c25gi/3Su8wHCssIG5JUPZJj9j5rl6D1feFp1lAIw3wr74sf2RscvYEGVea159W+
xSlVblBmB6MRdQVdvDVvwlmTfC3I755rTig/KCigygWlO56iyPzAygfTMUQ9OQzp
BvUlgbssbzKsvF7xjwVOWM9n50DG+XpR4pGbHWFoaFPETIpAD67R7xyb4CLmIa8v
ba4vVJ0mkmMgd4NF7+rvhruQ2kjnW0251CevB0vfB+D4Z9CiYbAUYMA97koODPSK
TDhV5DTolcYvxXCwTMilsWJM8KoKK35iXHuOecxzJgP7UxXjZ0pZGRSVDIu6x0xr
q25rMUt4jKkYZXlgMlBrQ+hxYAM1UNlolMiu2sdkVJk4ubT3JyYOFK6ve7+nMZjK
F5oqAOWYbvcQTVqUIOBaLCjgDOssB7GAUkg4yOJylUocvFOHzNsKQx3E+GMn/9XY
RljjDKWeyN+Ya2GpdqGPVBRjJdTZyCIptp80pax/tUt+m5v1u9SCF+9jyaFk6p9G
eu6LXPnuBgsh8YVj0mjaAaddc/jbxotqT8u0nCmJpibyTl24UHC8oQ97Zk7XmKgh
z9mcspHjN2saZWxjjvOP7aRANx/IUVm1Bh/AioKECCQuzZE98RtrQvTRQS2BJYGK
YhDU/thS07y75z+a5/TG7r0EwsB9K661QSRu7slbWlHzJBDnv77CgV3xMMesU0eA
dWQWstEJ5Gt/3NE6tiza4g10ANQ6bEEwbp6Mbbc32XgxdHmMX9tTTgM5xGRc3B46
5Y8gqGX2B/gaTwAsB8X4nnOVhLZ+l70vkUUMLCIYMu5AAQQZNYI3E7lKF904wykA
njEzmWkcVxNLoWrbIXhRpUhsVfVTTJBwIEGayz690yBiOSeMVlcinX7p7+mTb/1z
gmW6q2q1CAkZWIoH6C+AE75BuJ7Q0/dZ0b/i4fCXkj1YMlEYSNOCoSAD065aJe+Q
+3B1vdANxzCf3k3MywdHRz9JELsfU6WQLCrk7VpsNqiixBnkSbrmtS2zMyoXijkO
D8M4Rc8TEnYfxDrSGxWA92vSDRttu9dXjbgBm5JVwnp2yLyo9eJHuAwPJU+oB+oH
kFbot0qowFqrDz8n/LsYZ6mXYv86duxs/+/Qo3hs0cYRqFCNrUomxOSSOJB8KI/0
/lk41OL634SKuS3zpgVrMmSMbyhVAb1pDVod4DAr0cquL8NDAINmnnm0bf++zau2
E+IIE1q6GUjTOcfKtniUy5AQCrR5l6O9+Ix17fdOKGrfnSCIUFdN1XHcvfY8oGco
YjaMIgvuO951ZknHR+3+l3Ar+d+Ah+24QZYMgi5hgE03xMLHneBRQv+GOUB2bI3w
u2io6xwucm3P54e578RxGwwGqvh+Fukw9R/YdNmv6U3sDk9MVA9TzTnVGO3bfMiR
xZ68CBeqVaft9qoJfCWBGjqvCO4JK04eFMECWK1swt4lkTE3rQsu2NHZN7fQMDvJ
/3d3OorqSAEtBjwBBtDfz9AunuhmMN3ioHa3ZHdVprALV+zWEMGZmDAMgoWNVAqZ
Ew3mdq1oq909Tm0tjN/c2rQS/HEvg7u/NSHJhJlPfSj/S9s2VoiygQWjcepOyfUE
M0H19C6KXkmzCE+XXXPyWI/997CdZ0anYWzEmQiU6+8r3QTcm3Q4zc9LHYVtReix
CETlzXEpbeNbJAUHgSbssolxsDbhvCWD4WKkze9EwkvLTwGy1dg29YuGGIWPAa/x
u/9hoUyaptvcN7TXyBUh0aJJhTS3PQyX28Savixk3Q2g3n+STYIRSesd03nCuPEk
r+c9YLmIWJz850uggpK3wTBAohIt/Inw9ZneXBZkw3tnNWhIKPUXmaldvjL23OOp
FGtTMAnhR4bSzd608r0RpKnhze7vVZHXtobZCHdgV8PEixkjaXlcXtzBf8l3Zi6n
CViDsQX1S0ddI3EZ3wAWEXNJjlJ8PO1p+5PQhRNOg6pmgGJ1FBjwHvSlVudNDr2j
iZy9yjg6a0sUKVFkIa3Y0oxQfSOXBuoBrj9PK9MmB/9a49tJGAsZpWvp1+9JftWg
rT9SDwSX6TA7/ELNeDE7GRZMpHt2qo+IpSfOJUv4SctE4qaTzgb6u6b2jje97DTj
hGGlMacLu8tYDuUHuPtDsXt+ALyav+YbZHAgB9XLdqB09ldUgSwFiaRdNJpPWGcT
EC6LBVrUTAjHPSS5H/vYfgG0mO8Nc92Sk54SplYw7ZsHgOBBLv1ItQnwRYCXk1Yy
4Am9ySDwCCq6RDlTXsAqJLrViDt6Ev5BgaWt51EJT3sWUVrt1k/h1KVNKNaJsQS+
aIP5MoDYi3iVNOYduRYxWsB+8cOhQXYeVe+HNyQcxngpJFAkdhBeoSxqOvgTCK62
nTNt4rRyHAsXuzbMRf2uQfggdZ8u7BFE32Ibodxgb97wkDKK1Vt04+kQOK22vzbA
IZS2XvQ2yh6BZLEL8GTVdgFBnd1SnnFbYWCK8bnZNDwzUPw4UMpqFaydFK2XOFl/
Ibb9sf//gv5DlOEYOmKtIYvZaA34XTD37pPHWIhBadsbGmic3ng5LMaTRvdw4YV/
Fh4XHfKspm8wPuk7/hkEZUf/FC5PbU9A0ab/OmfBCgpzsxCrYoC2kKp/Uu8yBIMB
tZnxltjVtXiXXrEkW2tS6Eb4K7YNY3fGPVb1d4b6yQqBX8vX9YeId3V9DM/s2jZG
WLEs+bRJrW1Ua4PJUwlJMnXW/00mE4R6AdQHU1JxO4HCjsgz0K9WFRitCJAgxPPJ
eUhet3QIlPq9fxyf93IU8nwoOinAjK16GcfD4y/Dc/O42w4xIhU2cGNq7dVj4rzO
QNJboSOkX/SBuIDcWQwSVhGhRcfpmnWQSmBFK6OxHgJLuQ0/FC6o2a2c7b3pxNjw
VkFKbEKzODrrLSmeFCsIqj9ZxtI9eDxROi1CAFs2cFUzkBXGMFX+51sVvg2b252x
iqkhu7eOnCJ2PmEIZjALRkwR3KXkmxltyUeFqUJbmzFyV8AHWpV3WKneOuIS2Poc
urqTWgHI8S3YcJ7s/qDW9/96Pv9T/QS8N8RKH1OB8QQUFwRei6WEIk1EcdpDiR1a
6YM0bfgp177Zxth4d+qrVMNQxBkv0/bR91caxjFdmJakeH+STb6LP0f4WlKSHTsI
lrhtRnUtJ8Jt8i4B87bDDG2/TrFZmBNG9RYj6GWQy3jxOyjBkF6Pt4BlY2/8gsQZ
IXaM3dna59IVgXF95JRh5cUKizNO7G8D+qbmZti5vO9rXOQDpOB7QbIL/n+lpKAy
QPQZiYxwLS8esEpbP7GyDqFueWDc3WS9L9XZmRvFigNYS7V27qvyQNbFbqdDrfdl
O2u7oTaIG1nqsdNd2L2tr3MNBzOXOr1WJHaz0GtTGyzXgzbBlwaZZK+y28d0bf49
KqVFUR4cglN8WFT2lSKa9bYoGeOwy/swAfRx1CPqW2Mvw2qj1rxZwE6k+LhQxwcw
FNXs08C7XiicAHM+xYGIxj5eNDiHA9+Jcjw4wZI3n2wxtYmx4G+8lmuNjw7w4Px3
epWrTFKdbxKkPQzPGCdww5PcVOcNsWvtMUyZ4oh/rfq9UZXDOZaYs9C2kmeMhWH7
yDE8WqqSvSVexyJwcKyspCepIqIbIQ9YirzTp4N6gsTCidf3PicLtU4FwcN9tKIg
KfesrxpzDoi4DtF4XniowyJSDa5IvIWvF5kabLFicIwzaKXZ5a1S0BqF2ey1qhy9
f3vr1lR6Ifoc18sDeH9luiBWuedWAyEgnAqtHtvOx2Kmcg9B5L0NK6anpZLq604H
fUbtoMtJ9g+t7QN0bcTQU87Am9ysLO/Kq7PhURdJ3/C3IO/fD4qNaoFvzyoZ+DVE
IlyWb3N8+D5VPdaGTafGlsyFpNIXuquKAV4O3J6Nq04R0WBvKwQH+S4x8NEMIIhf
VoR+SjklAQWmzForkHT2GYzBE3bnJ7Q+stAbeofvYHtOEwtlKPTOGa4GY99mpPat
Jn3ulDK/D2p40nYs/Y/+JXiOV93VYDXxGtEe0uxxN9JFe+T9MCuk/vaivIDXtgwi
Bcb1zFdn4Ka+5efrKwEnWgbqHjbG4qD33FMQ47E/htCmUPzTIjG1Z6/wvWdSSZDU
xdZWLJdzyIwidVIHsq3Aln3z9me7vF4zM66wWTuSVuAVxcMHAA4850onOtCd34BX
TzQzSSDSZ+eaUJeTPNz9bh3BIk8Z77Ho1M4Zl9/PLuNnBcOKlPxjbPrUaaQZK+R/
anJj32T0slLgQJGngK8wJTgl5WdJXoF9dOcWi+ZRhMZOYJmfTzHNARkuYJuU2LSO
JpVqQtUbBKbM6oi0MEIVkZ1XpOrkiG0j+d17o+L238+EYzrA1HtWS1Gjdwc8MhD2
6VBtHGf0KlcO+KF2H+uosRzDBz11IM5IONQdNGZaydp/RCNzDWFab1hFKhnZWRB4
JimYWfzCFu3DmWaANqJWs/uZ1d1SjfVFL6eWwEewHPLUPxRjzcDRMpKA/B5Lmit7
Q/DhmdQc7J4qgtcT04YiI5CfAaA8znKtOujybo2CnySdggcnB+HbSeGvgtTUQx5h
ORzAMBlS1JTW9MPVMt9ChrzwXbfz76Unha7/bRthJ0HbD1v5dpA/tCSg0uQ6UocW
Nwf791gZ22YyQNczjTDib4A9vw4wwYMBrWGmVgavLr4BlnsBIpfa1vjVALX+PBBo
edSTl0ZhhmbQqlk/3J6hOwcBXbGo9kHYLdhBu+Jh4tCPJ+HYDuDHz+vhJmjQQQbd
NHmHuen9jcuEb5iSc+22smAVU2Yoxp+EVdA4Pez4+vdpg9F9F0nFOeoJVY4/AiyF
PRv8N7G92N54FTLf5rrHXUkOXtKY4gRx8uiyGsPr7FjyqqLmkciHcybj3kYt5wap
ABlpfgeXTsAhJKwDtIxcGDjpxD3TLwTF3S91SxFgv5ue9GunCyGBCVRv0wl6hf4i
EW5PY8VABy1MUI6CmRN71SgDX18ccUUSCYMf3hQt/3mwxlNeACfnuAWOfQXEp7GL
xXPk5ikrSTWTE9ms7CR7+4LPaiboXZvOGZo2KVc12Vau9QTAqpaQv00uIQbcHigr
73/hIzJLjzMHHiYhCvG4y+HNk+Y3R52s8iZuSTJoEK8ZhxYlfJMF4lEwfSdpZZBm
IrzybASHnnUPl5NQz0z2zRiJHmT/UKNFg6mpqDTSOKvmjg4aAleGC1zJgeb8g7wS
MygEJIn42U5afFlLCdyWlcJGAqzI9arVh584qohLaKiD7xlKVWev0mZI0JaegfdP
pVMgWG0V2d0UbhZpfvjgFC4qXA0MsbUvM/JOH/pJoBPFjHaUIc/qHT/iRYULSprB
ePKShVajIf6+fc0UzPqXU/Ur2QEFb93KFEDLP+pDGzKt9lDoYXRvLYfWeFZwl2HK
9sQfnPKGF0vo4gt8enZ6blDHOzkAtp0TmZyv9KgEcCqBivi9nI+0LgP0NkGky3Z/
0pdvOGL8CpaU0wOSwKARAoWqSxzLh+0i7XL7qXW/+m8YRU7DXQ+5Vv6eBAm0U4JD
EsvdalNHyfhKfDMtXNS7jnG9THUcnxcHC/qO29ZpLWinPmjNr00XvdvOb4TI/u3R
H7fK7zosS46LJWMRVHZwcffe+gwTEhCoYWKMI7IqIZYHwIC3rs0rL3klQCgHXl4v
QgcFY0zX9F7B0wOZLTOAt42ETqObW0d5VpV9aEzsP7Cyku/ZJlihXMQi8akHzLff
T4weD++y0mt8skqnAmyYS/hxfVJyleB+G5yIPB3D36gYpDXsl5+Otgn/vLKhlU0v
6pEHO61zKl8VSneNXxIO2EA01cdkAwEX533Uks+yT1exG83rJzSgADx9/XBZiHkl
vxIwwjHhBdbkTnKJ6hIRCIE0SiIxcLnf8DINvJVajTy1ur2n5TOUnkMfoeXoRD4d
WnC1Pj9IYUbN3KdOXsmq39px1+3tMlHFTPDDX2iLKbXAAHv9+ZGefmDcNrSoGU38
O4YmGgzihKXLx+XhDxYL0s2J6FqZKUFw3nw+h9p+noLVnxNYnjlnget3eK8k9X+S
+hndX89k0lW3lt/NoY3bReyjFzbqM01wRgxqRtbiNuJIDE9Bsbsp/79S+/ClCsGL
VRSBXbMDtIWxSTcPIqePmTgJVS/oEICqPwWh32zWuMIDadN6BnKX8Bthv45mHSvn
09Xn9uTUkFRR4kiMCWhfH5rvKU8lXIN/RQC6kA2g1ChOu6edTnkLeuKBEfRdbTMi
QbdtJaTmrx6NdazwZ4kRW2fuXRC+wsdedSJcWa5ZKIZVaB2bvdTIjqGFvvNHtRtn
CcyhO3lSY9aYJ3LKgFsfLSV+xWIw//BVCW003tYhL6MdS7UX4yHNzi9Sl0/DkXNu
qjv7Re4MXQHIhrOQWDxac4mJetZCKANiv+I2PM/hMRaPtkAeeq5f0Zv1IFpJjGH9
9HD1xZkzUsjM4mp+BIsfbtuQi+nwViyfko5wzsiWKPNMtftqpymBu5PBUwii5xzo
rRg82i6tBCpKmqrDHrFnRjxHZwkIMAVsLNqgpt7rseb/CdlUd/S0FzYWoQOjbqgR
aEoXkVcPlQCSKOem9R1iTrb7Lbp6jJmFteLEQMs5W8g1pTDA40BxMLu2wartLNl8
9pKfQwdIn8aDCPXUfv4srteCftsrCaISiJJgtdO02JZv7dwuySX89T2J63DG5WW6
TI8gmB5FZMgikH2j1Cp1fzQNpis5cImqyllB6s8TtyoryBvvcMkeux++mQ7sDxRc
veaN7XBLqo5rPSl/xXRI2HZLVqW+cTwaLPR/wXnVpL0v8BVUKwtgU5TrAJdeBIgQ
lKJYVKTXguFYFbP4TZZmvYAybzUszCTNrbQ84piz4ULnukBsrYor7+HLmo53Y8Bq
eru3J/U9oi1O7364fRpGgioBcEEZ1Spk62v0iFmTNsrgxWF8UsUz0D27w3tbU8gg
plQmBOwm3ud7iXRn4lDVGDWsJnOodtUqi2T2S6MvM7HoLGD43aae6xrzT8SWiBiJ
LgW40US9YLTx7NZUenQRJJP4l+hYLvzQ0aavuft0Vosccb9CpYsaV1abM9JJBQQr
xkcx1uQ1F8nP1WQ24V5upOiXfjPegqAbOmL2SJvtZ6LniRj9PxEe5DbQcgKJCbhT
gO0QDyr1iW/GaSh24IsWhVZk3+ym/T9V5Y4VqnntB+Pfbo5qI6TCzKKu/xWKjfED
fG26VYf+3V7bdFqwKAbWc93yOKsjcp2lGNmLXKyf+vXTw8Re2coJlaCrrbliqoie
BrO8B5y96tGhyVGevpbc7ZUWoJYqbQGs6ySilJmp0gCZm3UwFkiQdQONc72YgrPi
L2LhwlgFJAltavpY2cWJh2NaEzm+XNgOfNnAgzaLtPMRPJf9dbuQUz8CD0HP0uJl
L51QjTutfP54axGJd5aoCMffQWz9cbsQqG+FnKSoV8y+8LkxTkc+maxdFA6xkBq5
MBMmm00qmwrTfIwFOLlta6DWe2yYuIQOEPoq+OjtbFsmiuLchBy+btyfkhO5s4qh
a4r7m0rIHPO7bMkaw8zcVMRltaaZhMeu15CWZ5JRD9HBoNogmS8lJKO91Kr1xme7
Dgx6CKlzCFWV4cT1K+yMBzXlV+eVggm4RIKDzEPK6LKoVTXkeA95pY48VVD0c54q
BWTzNyDQ9mwt1I4guak0FFk3u2eOqg7xgEzYjk3tU1Bo6+4LvJKMbW6iIsY4Nxl9
Yi8JS1jcZvxcNcTq40l2aTAqbTdVrqt1ViUmwUfUBvRz3J23VsT5p96R0blk9MQZ
f6zvndiTc01D8Hdi0SOBePXDPasqU1uzF4D1pkicGqhWggX1e9Dkq8kFE80cx2sp
uvZ7kKFpZakBwkZ7cyUOQUzQydFpIRSSHNyT6sPspKU3g/pl9ZTpA4HndMVQdAya
WrXgwg732ypSPGL4eeNsQocqvC75LPDK5lPysFSxBi1Dk+jxQDCf3w7Yfhst8FWp
idwsW8ZAoZeipUhYfcM5bGVunnK0JtAZQFrpMyQ4fZ3bNASktPPNaBeMgxakQtIh
zBTb7dx1Spn+hmhc4CHvAhVLu4zSEhSeIdxPdcAzact9KLiQ7MxD4l4Pmc1aH4iD
CljsW5CAs6zn7kmeL6iR2rn6BHTYYn6FQE5t4HNnqLMxbyKUa+nvHNcKqRY8vJvz
1K84HrzH2AGwQeqQBeEXVAYDAUvoPLjZlcmjFP8nqEbjUMRt5+GutAvSt/7SiFtB
NQ/Vss1GdQ3EBXiTiTI52Hn0DewtIvRz4gBU/NQIJ93psk8PkfnN8LTVVAtenmXV
+Wq9dx+zSFsxQo2FioMDFXnyXlTTYwxdPJ8brHPI4ZzJ5/37a3Re6msNQzwHRP8y
UvjJ/wOEbFsxiO6ye6ZVTCGEbZswISG+TgjbruY8/F73PHXwLt+w7ni6+2OTnCK5
frYUNC6apVybvfgTx05Q75MvZgbT1v25ZWVEL7H30de0BBpLQsrTxBMVCOo0gTLP
2ucYJIU+bODARYf6X9GEC05weXzhqYb75VoYw0FUP112jnAtoAka4V0siO/1VQke
PKpeqP2XjsIqZuDzz6DgJSwxXHNq9jUyxwB40ySwhubPjU9+pTRW9r1bv3sDLwkJ
2AbZj7ju2N/MBz1p4zFCYVxdc6LzMVRXlpZCx2hJxzNcz6oiBEA9XtoD9im8GO9Q
NyxQZINudJQvLKIzQdIL7jCHhHcKvVyrCusLVOR4Rn/tHvnn3fq5LzJoH9OD4mps
mP5suQv8UOT3/CxZ/cXDhmeailEZ6Ng9u9oE0rtG0bSpEVzQSXBqHavlmUygxkab
PS2wTW5HWY0fJ5d6cgh2Cf+Mvib1cRRkb7qW9+u/tP2bF6Qc1/Wgtrj7R7UJHB47
/Y5YwfCS/ZYzb1gXJRGrKMnyoY2oVyhK8+0rmBpOmsgal9K/Wgqq22FGEDUI3MK8
HvpS7HVsBm3xa4qM/pab14LkWMSmXpMe0IhjcFvefnY0h2xc9aVhrWPiTuNQ6d5b
7HB+EHSzjlI4sbv2K4uVAQjv3v+Wjj2c1MyIeHCs5aBYv4bjsF73ZQoCCiTruxNO
kIecVbMXjOjYcVMwDyBAwcOW/KMKPC3vENLwRTadi6WwW4/HE7/EzGEwvcNGBLpA
jvW1g2F4N2aRaBHVLyxVPuugnsYUX8d4YhbG+4GwSFkLgL31MALMoqztHWt1adBk
JTtIfcxC8XMSCeOXvFG1OVaXFsN4QU6uerUHFmHMsC1dhyKzi+8wgb0RhXJC31d6
idESMlwh1uZkdN9paarmQu+nlQQGUcFDv+ybF4LONaXhQ7uLpaKXtph7Yb3aCTdh
CzQs3x1l0YGcY2rR8Qge5nYVcQwdQzvOVBWQA6uOOCekIyyL3rUm3MTMhsaZauag
AnKyW72Md0SL/KRlx2rPRGKOCHUWBGyM8KCmL8suhye5f0g87l53TTjO+35jfJ7Y
FfDyWcbKDjb0UHUjIybmtSRW8BjiUbTxk9KMge3ny6tRJeUN98T0bW1SDdiVhJDO
ljhDx/foso7LYeAqvHYqmBzISjRrSsTg5DxU8o3K82MvRG0lI3y0BZhwtrTCeZg2
Vq5u8hP8rlUOUTV6mS4PuWP1uOi9xEXayLGw6lrmHbCIPIYvEx/LVEwPvpEITkKS
H59lesAEhUVaMv2tVsC6b4fI5uSjdwTup6XFufJcyqhhzXdKU3WLlhjQo2IJNLPJ
VObtc7uOodrY5qm5gipMFL7bcR9LkKoniTow4Ie6Na1IaKYykpOEx93S1rnUZ1gG
9pAAKYuoBCIwnCFiWZubT/xnaE7kkcnzHLxFi1D12sQ8Wxb4h+a1rnAga6Uzy8CY
UEZOUPCLnd8aZgtjbg2/i7fiko4ltDr5btK10b7R/NB5YVTZNK7tPyfg06Hv3ut/
ZVA/latEJIQXJzGycwY1V+tOlGb3BwVhGbNwVh7bMg4YAgcBkRKhCtMque+W/fd4
xC/XEtkbXwl4g6KRNZsw/FUnJz6tBfpagCt3f0pRyQ2waLsSV2QDwmRkJ+oMbpXG
p5kMFT2QAVyprc9zE3rdP9hbCbxOalP0vumq7r+oZdDRPmgXlkfRhnwPGFGFgzwA
0Wy4SFRXXzHh1Bb1Eq01kGCsYH9U/U7erOObnkyYNxH6gb1WEZoOpFwnUsRlUGBz
7BkitidIcqAcALTEOUt4G5WJmP1PF7+HcBEV56ExjlhphEpzY/AM+lVayWqx0iNW
dxfcJpea43ITaibR6dEUd2DjCpTXGaLqaQB63tOfn6ZmoglHVs+TV8EwCjeBluCr
m4YwRWJcZ9ZH6lXOW3wzfAVDh4Ea7GCwk2MX+JGgiQ2IRbF4nMOO9zmwrrV5LWO7
3B49CSuyj6/85auIfladaWJs9wneT3gjHOSYurQlzrVsF8y2wMt94OsDsNHJSPDM
yP0TqKtjqqfVdfKDSDsTbuoK5JfQGjVLymZvsfqalp34KQDUG1ltYmc1q/WZy1D6
QiwFzvA37k6tFLp+aJPgARf1HukgU5zQGrVRa06yv9BFaSJe/N8QIA7Aq45yIbxA
E/4He9puaI6/UlBcw1HThiawq5Lg9lZeS2klRPyb4q7/4GkAhIQgftAyAaQZ9RRP
0jcaut99fCrdEEAs471iO0mNqQ5n/nBiBd0kGSJ8/E/I4xqPRSoVgFNvKwroOZmc
ZKea5OtFu+4f58nce2JA/TAZQdVFpISn+X+5QHuHuhizrM/hBDmAgNOnAOj/Ay1o
UR6ecGHdRx/nCqvsB0rGW5+soF509RnNschZOOCcJx6iR3Sx5/6675lopVBRqC0u
2eOR4UMMsRtkoEhwJjMQ5FvAooj26Np2VL4bfnTOvHG2TxnGK4YGZYfEMah82sJF
cjd2RxmK8DBic5tIn7z8PbKadwc1TizKCf2zbr5clL1160cPF5iLTIXO3Cz63VVz
HnOHdXzdqxX8SiXHlgfYYk0dqoxgK2KlxUAI+N58Gmk02oMVujpWBhr+ae+/wY6y
86kxN9Utl0hhTmKdSw3AYiIT81xFj9IduGpQLpDdHtUd2WOAHSzrOBgf00HCqceL
m3hrvoT01bL2KtZuZx9zENGd/SjtACsyO7jEv8vAyYVYiOV0EL733EcyYs0N/Vd4
X/SD94MNTdv0EGr74dTwavlToEFG7BBXcA8/mGS5ZOx9pGIsf/VSxGzNuq/dHQjC
IueluI6bHerpriLaPfFfz1QXVwNglRRwnlrZ/U5S6YfIKUj3Q/eV6D+sAYoHZhBz
ffdOdBZ3jpm3PJRbJf65VSubwO+awSyuPFCHW4wMnmnfllNpV4wY1QRT5bN/0qQX
u1yHl9XvX+nTWlz3cWBY5AaKFDKj+OXu9A3eJBEFL24u3sL2TcNHN5nzO5PTjjWp
yNfepRXCCeoOPOgwB2GHiRTovjYc3HLryexwj9y0yC1iAO0/VarAad9lAx4uN0BI
2YvsBrHYsnBkpQMZA0nyX2Vu45CxahD716KzNuzEM25dqtk0i3s3MdewZmPq/ptI
u3WBXoCIqW3H+XyuDbXS7eEu5eh4YNKlcbW3Qo5DmDkDtTcf/Kd8QInguDs1GlLL
7OmQ3oCM4551tZxSS/NxQitqqUcEWtdNw7IKMfvZ2ari6uNs6OsQJQrhXaBR8jYi
depgBySg0horYRK7tOj0N3CaeSOIwa1n55ShSpkneCpiTCSciB8AHluuLM/6yZbD
Xz3BaRm8a1ADAEiM1VBeJ2ub7+D53kbhAYvtNjd/PNno4UyGoxpzDrPwfkHeFAok
q5jWicRdx83AQzIVZ+I8uw+rqHip/LuDPnsXbD9J9I+gDfUO0VLR/gWU601MvPT8
XgwHcx93zXOVZhRKVIG0eRs8GP86D1YNAFH8mVj9geC98sw9jyFqCPHAWL9SD384
pIYJQF8F6BSYzBWIg0D3gDgqZEYS5K76xigVXEu6gMAMS35U5rRU9pWlgMQw/EYT
FFZLz6Qfyl4y3MKWKToQNQ86BU1AHzvyK+9/uQblOGXKtrNZRXqZ7kUoTG3z2s7T
RzjIHJj4n/WPpWoTDkVFVTkRFd0/IEyxkbMIKCqE/7u8Ss2xPTz3Mrhb9JRKgD8y
OHXrdZBs8OlrkU1vh4jq+R+Hcnqj9RHUX/nVrkYEUenidDzhklhIHHInXJeOvlHg
eM7O9Idhbyok3k50D6SXZVAiN6GW4nAQRdVuU/rR628Iyj0sd2qlUPQoP8IT3z6C
Er2GU5zHcCiggKV5wvEQ7Ny+bVKrNluu6R/dxGT7BM/cmkVYNZs9ndx2Mw9pop73
o4Yz1/05Qn6stU58ROF5dFVTcoC8L7TwbFzi5POl4HJLfJiNodRORi0RPLS90q8k
P4af2Obxxae0VFKh65SWRDzKLc6iauoeQ36IOU5k38qZ6or9EJZex0/9Lr1Awe58
Vp0dmEiVGMsf74J/FZ1WtD3A3ZA/2ImJy9VE0U36MpQmwh8eQVZ7VA/xIxwr3/kb
TXtsnl+UCto4GhOLNXh7N07pRbArDcfgtP83mXDonuLZD0zqMEdlg28dUnaVNwCZ
sbYBQ4oftGFZ/E0+8N2Y1tFyqJU/3MiUHQ7uxMMchSU19EHTRrGScD6sPFa8vFPn
wle24wI9Z8uBggkAHMSn3Vy2Qt44kuh7i7hN1QAKxIHePyIZSbJraMU3vyE0OVd+
baimf95fZEohIUsdbWbBX0rsT6styX7wrtLRJhqFB1ZnUVd87qO1Es/yQhgYojQV
MYtHl1hOKiaV44OCw7I5aiHVqchqmsMfZZYCkeOLBZuUFb8UxmQXBBsbcAOfuNZ3
yA3/yqUjqqINq3JveoQjVvrrhaESpFMicOcQ0oS02SyDEQTnSi0HGcd83FuMeQVH
BmVIpHxT7SLjLqR62T2GuZXOYe7+H85bTqRMOF4jN9KDQ2MbnEAacdFCDptX/1Gq
URaL+YwnRKlSLB5J/aUKg6CP228j8KfDEbbW5UkCo2OxugXv74rHQneC1wrL9Gzw
aaSQJdAtZKd7MHlvXM1jJ3BdTMql8/AOc6i9H4Ra9u8SVSmdd0fme30QCL3NP7/Y
CxQv10uDX6YU8xWtGE2t4RqJda+SCcIJKg07RQN4OL+KoeZy0KV6zuVN72iVdPSV
H7wd+Gg6ReAOrj9RhtT8kLfR8oqbPjaB9PHpZsUOriZDlTQJPqrPZ6Vc2mkQDq3F
eXPR6fRlGsnnyqKoBfM0rlI1uymj+tMMuV6bsE+LOMwu3AdrwPHeg7fDqjYX8cpx
Ga3nPEKDyf1+0SqvAnuLSqK5XACjLElVpFRgSe1CzMmgp5LodQkyXX4kDaHpHMr7
cPN4ZSLua/zjX6Mxqy3lVBs0qoOx7IOCflt58vWpWvPcu6EtftzmgnM/adsJBNRr
LRZJpymL1cZXf3yfeJ8f6to4ybWU6ZXkRYIY8vIfI9TwVtplxfXl01N0E4mmVsCV
y8Kk8xALj5zRJ4BqBbtS7f2YzyqdhEhSBVrkOGstIr8+fsECmE1/3REwJURO6JFk
UxYDAoFdDD7WNbuMMhBuYovJVmzlycYggX6hDRSmWpvx8QbS4rwYrtBsJigFq0Gk
x/mhFvhO73odkqcObrSkgpKX361xdtCEV144Eq6ObNXhxI5/5BVYAEDjmoOSzrJE
Mm61SkjAN6B76flLelDKiOKtRQyqCcpYuVVPu2FMPYiNhaIzzDtPaI2cyCKxilck
EMsVmwDIqVLiUo1UwBfYpnS8gGBYag8HeJxn4WjQJMbNZo4XsfxHaCS2TXXKi9Ex
Q250yNoXLp8WKdVKIHa8UtSuoy+RnuNmhPq343WwfUJBNa7LXwzGCfTf1wt1wJTC
mEWlK4czelFCNMO6op5A2iGuZkfNjz1gN47SptGJxvlexO7KPnqjZS50+3Yu/2y0
FDLeZ4YeQDfgZTL+WB5k76VHmFcAVSug0RsRLELGwh/zHpScx/SN8pmlYpSR5wf8
gFj0oxFy2jcs2A5KMH+q8uC+2FAbN9FFBow9eaXu//RkhRqzTpS4PI4TAax5LVae
EJyA+KxSRyHk9KU7fYg8ZNXf5hvNlxevW7D6R/maTDX7/23NSRcDTEOKEdkHPA4f
fosdi0eMx8CVpExdn5xrjylCMOv9clGVuyrUgwm9cmvYIC4m+c8QEV8DHd1+MdNt
6vlD5JBRzFsknM4eft6AFRXGx22r3/zijLN1WH/TmJm+AY1dpsKx9RbphST73On9
nlhp3hg/RgfvltzljgE3oaJh6+AZstwORU6v0W4qoPJMs3Lz/LmPl2rHpnPI9VCe
vzvHroDKc/ltVIAm4t/GdFf/wo7bceAWKkPn7+ghtqjSumUUIapLqmR6UQiT/Jid
h/351DywK8XhjVZOvvFRzVAaOz1CiPTzj5DR2hp8fNqBe6bsQze9T+nLKtjkQBB5
avkZYxscbAkjaXGZA3aJQXcQzYJX2Y//KvAPTeA+0TnO42Slv5DYZ8K9UMVtLOf4
xGbLNQo592+N0NULPq41P6NQ5ao2LnPRzGXajq4toav+niZsS+9D+fni4I33cQCy
oN4TlWrB4be8j9gAq1WYF24K18kw5BBQDP5rablJTNWXRUe2Pu7gC4+3j5yr9r/L
Zvv9SuwzpfdM74jldl9qoxZ5oS0A80g10y3gc+XeyWCZsBKTxlpsUHDitPu2TGEc
hj2oypvG4DlTSU/cb389pZLbKJ7ZFkqBP2y974L5C8UgbwDwNrNsX/tUILC+ICx8
3KSq6yrd/GJCW1wqHdT322oneQwhiMH17VqFkD3Bk2fw7gEGBJMm9GdjojD8RfzW
R5xNeDo8ANe215neaIOEdN25YOJiwj49s3UUeO8ZALoF7HMhT74YlOqhmY/C4w7G
Br05i8WUxUvR7v6g1jS/L6hVScKF06qpZ49OteN01TOV10MQ5uS7ua1Ma8Eb8dI9
atTc+kVSbTWOqaiI9jeboXaZeFAkN13OgiBIM21mWqLNaAIHfqADPCWIqV4sRUF5
E/PosnEzbtGn+BYzZjmMOJ2o6kLCpjrZaZ3EQbipASMyY2zoJQDT2U3b8wN/d2bv
bfQP2dQccrK5yp1bAlnuvPtNIuVR2NR+7fI3AlOip3jmLLjuKhb92ZJSVh2v79Gl
bCj8ADrIgQ9U9vQjfG2Gaph/PKY3aUn3HN0f9ICFwmntrrwb+ef9rAf3IR7ikQ96
OFQqKp78PsiWWIMMXutMWU4k4VpuFS217iK9TDmNpkHG0PZ6+9sw9zFT7DLmKOJC
JTpgfRq1GxvjBv/akqltuU+HRTDofyDa3RO6Mbqum1UNlJhb1Mt8ly9j7Koy25mt
qMdEr8pDqtG0yPcEswrBwr29frPO61p3Ibkp8Pe4FbTr7W4d8GIKsztOB1GWngMo
YLffpRp8rYNHqfINmx6ONoE/673cBmscSF9JoI/99O+jsueGrRPieL/ZTASt8x70
E+n8mCfYxq5HCBX0zr3pRhLh4pREEETEQjDy8te0i/Y+19+SuFe9nyCcHsa5mL5V
lBHb2Cde7N6FZ08sCkkkeLGxSsh72Gyeg1IUVxNWiZUPp0a6Z1mZY64y5LoKZV12
prDt+8cZxfdT804ZzB3xy+ZAljAJGaaHLkotms5j6eJjjJmby1XtwDxvb+0+LLEj
a/k4IjU/DVF4B+YFk1cg5PO+1JircI8F2py36YZINMYxKaq7nfUwV3XxOXBRhGUQ
OrAaAFMiFUQ793PjZCr5k6qiQEcmsRlhsJa+zLXBrIgioOQfUz234MgPveF07TJc
8PT+fKktEByEBH/G3/z4aG9Qy2XP4djh/73ZVDvbHngClA/i+hbLLEdBlV4KUEtI
UE9DGxygyutROmX6BzkJNIpAukX6qcUsebT63Rh8rFoiO4/OebaayJVBf5ODP6h9
v0EZ9YG9fclRT2mBfj4/F0CG1avX9GYt8KKz36vsmQ0s5ldspgQPjeMpjIPu4zjg
l2QSnCSalcdHbaBUZmNwfoG+3I0waLg59DlzjyTuFoZ8MltQkhfxXJuMs8DEvobn
qaQSfM0htbGQvkAi20tq7I6fYMCg9HqyWPRCSvk6Mxmh16U3riRJlCe0CPItx7BQ
tvsniNqBTAYSC/VM0DKFufAdobF6lEjzHSf5cW+i3sGjbKir/u2Mq9N2mcUjMPfg
56b9kSFVnZWC7lUzg+dUOrfkwdlC0zlDatH6yz8cuczAr6hKi7Tep/792sm7IhL0
f07KYaCtZHi+KenUU5PsKyETh0DxMKzj9tmEHzPL8T8cYd9BZRCpwpBFuri8urfH
jqPt5fNPEs/CyoDOT011F0x7/39m9rew6b2sDAbNW2ZSq5iKkxnnXcYKvBpKAJSu
9CD9ZLPE+1Y0BpdL7SsOnlYwwIdUJNqvKS+bWo2RQ1JoLYVZgFzw4nKGRl23AGJw
NveZu1XFxKYZ/VLH5vE3bHScf3UlGxytEVp1E0uph3FKM/OtnrVJP/M/LMsTBeGI
HikMiwoJpV7xCdsuiyD6Egm3Z5OzfiIj4ryQQzvchpn/JC9uCYFika51tWiJvrWP
ja87VLAzC3qoeuBdNRacPEDmxZHaBxjinWmMESQ3H8xZeRYcwwUmMVQxa6WEaLSZ
prte4wu/tF++agaMCe9E1SECNrzWYIauiMRb7WL6umcaGsbCo370Ixve+zZGtWR4
15Lvb7W/kelEN2Qq3z6SnNjKKz+wZRmiThOWRh6Wv+o7qvIebSLHeZK5EqLK2OpZ
8uDj0/qo5jM8y/l6TMP69/f4LaPegq5IN8efYouTZKEQNP1oOV8TvaNXB4R3w0n0
tk84pJ/d9oeJQEMy1scpeEBjZC0kX6s5HlqSb/cKrJo9WdKFoblsEpXKcRiqR0Sf
BNifCouinpYvKdM5PZmf4AkNEaEnGxLIbzAClOJhIl4EqoRvCOqMGjLkJB2l6xh3
2QCvclvNE8VBNF6j+iJl5GKE4gYrt6WGXmPbsoKB8Y4xE17k26pzFzu00/85httT
S6P4NKy9pceFShlfHLOc1PA2zkS5GKXPzzVsr0md7/Yf80c9+rzv+q7dI6GSwHbc
cpAKGDscSxV648jj4AyKQBRpRohZrpeGH4SqYaDIhet5VPOKvSY57UpHIiUY3U3Y
Q07LnmPXWPdbDzEZEhzdYjCkMsraVDtOrB62BLzdIse+yQ1XCbOioIpX4MBu8uZb
xefhl8ZE3xUo7SoD0T7IvSpbt6Cs9MHiHOlbWulCzLBmoOOdR9sMPTtMS/5HUZlX
dT3xCK7Q16Pat9A8Y42jJniPPAM6tfzIw/69hji8sjAtXnkAb5MedlBWxAlmv9tp
Cpw8UxlZUG4MVBNIHVnvFs4zY0voOhlIZ/5AHurgTKlOLaKEQ77ctsqHsTbz/2Qt
djB5++R75kO8nVpXZMIFHTno8lKOrx1I5ehf/8ELYo4c2+tlZKtEi6tRrv/xgKNF
5vkGLMcIKroH86IiutEriGCrgsg7aZ/Ymp9Phrk+Gyblw6egzNshVTOfOqfKDmzL
zyTCs5hXUIB5uJosmFJl+ycmOMOskY1cl/5qMId4dGiNEsmhTcTNCaORQlWQvqfd
hboyqJrzGsFLD1xBVSIoBs7Fu+rQAzn5sSBFw7Tz5Swz6tHaMnOZU+M1ijcDrwcZ
CKVbDyxhhnvoFZEWatXTpeSUQjFhAu9h62k9N6XM9zh0qqIShNxkRQNjx3UQJDYy
t+EKoOF9RQMJgGKOoWbYvXdUKpiHA+KSpca88hI/G/c6p67BaVYt6jt0dATmY7RC
4p+UK9y6ft7zcEthJUIWUpiwTkYYznwanXRBrphmVjWspJSqn+ZvCvlmh6atgahc
77NpyPzXUtg6A5GQLrV9/UTSBohzxd0V1Yu6yWjNId1nWkba+59vvM7RnpCPaBx7
pacvKaM5iLr1MysStEFMe9vOCg467JZ2XlzZiMJYtRluEZ+w/x5BT5flBCr5zYwY
OGPYU1McwEJnlJh0b1VB/BuaOCvkY4jTJBiqep0ODp72F/rh2/ifFdDqSVpF0W1d
Wx41oypsBgGDC0sdorzn+OQ5oOk5pbeqRrmGYo9b7QQFUdwD7yivL9jQZciAP6+e
NAulP3x8C1UTL6OrnamM0FcwhHSVYnR6WE9xNApp7VdmWHp3plLIviKIWvn1kQAV
5okJINJ9xkL4wiJBZG4c4Uz5IZEMQ0o7wj34PgeDceMpfgJgD2Pne94Xh6Def+2V
zjbRXYfAwArLymzWPAqsZOYnrW01Bn3qbvs/wLgYwzB671pifJysQzQbgIobAkR0
nTfV05Ja9jajXV065paMTX5JNKNkrPpQdt2o/LRjS994iVSrn2srfQ92SrEI/9AN
w8AH0TycJ90b+eICAvq+KT/4nd3+vAM7XJc9crKT+jXAQwl13NA6CBazpcl7wDc0
kW7+4irELx6+spQz32pWhBvk9GfBrCIS4FiKCQ84ptSrX42yEz5tG/BdDr6QVBjH
GyfYY5kP7olc0TdpJ6G4UTcImI95Y9zVdhEe9npzRv2bW3P9FWh9do0bvuaOnu4l
1MvRbzzP9AEHQRu+l0yAeGAbUkOXyw1M7Mbz3lHFwNEh72KkWBkWYzpL+PC+ad+M
Bll6MvlRKEnnS5QozKc9772VDWEw1QYos+R9jIiX/RoNnR8w5o0XKxdp+rAyrgNY
v8ikOU0oUk9t+lExz0+1lZLu2M0L6CX2WFgmyMqIMggWKBm62ForAHP/LjQqeKdV
EU2lsrfcWQSO37KUelfYDMFL7Nf/5qDcBXGg72Kx/1/lOr3JekIJe/+7UOQ7dLpa
Sx/34Oy2Q4oQMZ3Z73z6LptAZV0TX7DvsJ1Id5D8ocgXtnrDbnqwJwHiYnONSdkO
O2GLU+ABxoy2vmFCuLpGAcmt9uTaWJbVf/HJ3N2cATxf4dz1s8ibQlFZZcxVwj6x
RW6q61t4F7d8GT/bxETbr615Zeeba+IMA4W/CY46uwhwsl6Uc4i9Gqg1uICmJiUn
0jyRsUQvaIOGhyoNKsI2lp8J8mQM5dm7ggpsbKwuWvtsQM5+kdbCSMKtnl5CD00e
1X4akJq/o7HyTXeZnnd5TjMhNPxlLvPXXRiEtZX/HiWZzZR7tSawEJVEkLTpdhqK
nnw9oS+NU0pAkm1li9+m+4LkuOrZ6q9WQBvokwVOlEgSp0DhQorq+++/Mhx29OJd
FnMN5cz+v4mp6PvgH409p8wE0n/Heb8v92upTzwmM0agozZ7fw6VUwQCElzgGX4b
L8NHJuZBORJGT0YLuhS3bTBqE2dmDT0a4PzA6VH56fnQ4NRuSnhW1PHfpUtf3SdW
Ug9325SamIgRl//P0HcDhwPS1BGa8M6q8FtYBHgrSwpMRlDgkz1LI41xqzphMSdD
dhCdw9+3soUv8VpuxXVCS8UfkBYfvbsKN8XIXWeY+WrZdJDZYesh/Q8YOgK8Fok9
U8bRVDz0nPQig5C4/BK4xTTeHn1noLGcI/x1VpeiD3UiHgvJPupVTAN73xD4qsIX
BOpmFVKit76RVgeE5Vt/JfqOIsVmDKS7FoCLuTrlEdpERnC+3rGU8+bAubxv9kyp
/P1N5ggls+xfy1R5g4+J+RL/UX6vkZmWCah3qClAa3+FSn4rE1dkCJ3/3W5llrND
wnuh31xM6onmSFmQKJu6EB/JMQBzMOrfLdE7rXI27NsK6RhO9aKqP/CM82c27SgM
XjOsRrmFQ6RXuXn0vfDHgGnCGIR4OTLVgdzIRMv4VxCC2x89ypypzL9Qs/cdQpI4
waH03WSmJyhNlFtgdWwxgWFjbfMXdUAtIjxnhEagD3OOvXxC4Fexf4IgDOnmkYPL
e2W58HjBrU9TysNHmMtLd7A0kvSOAbP7ykNkfOETU2teTaTEEpoG1BWPhSBQGtY4
62kBa9Q1/w0B/d5t0hiVi8NqxQf1WX0B9pFDB7Ms3Z4O4Osx4kOLWU1GKqg+DJJw
GCdxKTkIN16UN48HnleemijRY/CEG6acQwQ3WBYU4DswavhlGLr3eOO8JhvDmEwm
brpzHY2YlsIFg1pN2ohjLA29CF+qKNYWkD//OimS4Nwx7+wcjN/0iqm9M0pVaAmj
JmE5GuEIpnqx3g7qfbQlteYxDc5Ky7D7/QA4zEV/Obm/c9+fSIUUUcr8rGi5ZxWq
KQ8nzyXpfNCHt44fxCLBkcWV7TyJ1URr0jUI5gp3QuffFoaYIGJ6FnDMPmJw+j/2
/ZpF2vIeIss3FyElVauDVZrNUG2YRE3/Ow6RU0rqo3RhfB9nXZTeZw3/4JT6rGk/
OnY7roHMnypA0Od94Z+lANo1g2u2tkoAvUTIVkCUpBt0Gk3a9aVQbziaN+0bizXZ
qxyCQ3GFu+WghsbANwVI3pcrQSBVuqdUH/8naAlx/h1vxII7oSy6Dg2O1Gphp2ix
8SCipSpifG7i3mnEr8otsxEoNjGZ4tiL0bLrks2n3SPN8dXwV+IH1qHvj0JbPxHX
cgkII9y2jxJoEcbJCEcMbXfN0USYq0ee2g6Lq73ZI+tKmOp/8664U2j6iB9m+gpX
BiZLiu4SWYWct65R5gUiwo3WekOcscwmgXdRCtz5t0Iz0St4QG5pMkvuABXZpY2/
H2121DxCUSBiYCIsm4QJsYHWGa/F7Zs/9fP8PE3FiQ7Nck9EFEl6UzPKNTsjfB2z
2v+QJ+3DhM/taZMeDgzupOSke1Rj3XyRiMoZXsCBVlJgaGU0YMazCvLj3AcrfE4n
OFpinEF2tP1MeX0QnDZnUdVuEuNoTB2SxHdvn48yUXunpfZGhHLEX1PuQ5TZ02bs
7ZcTwOAdbHnx45UrKWU0n0mH1OArUz2WBabMI8ciZOeJ9FvXc+N6NVntHQf8ZMQT
hUQ9UDsRXtFISx1ARcTEDRBVrswOFxMC4+YKLr54EImNuOCbPRD1RZ8X7LD4xX1Q
LX3v8oGi5yQO4qC5rjvMxqZEZy6KvwYX32dCh1qnVp//1M3wQiD38+d1RuI2MrQl
vNML1og7H++6tJAN/LQULkl0VeLw5ODaWZ9tWMA2b4WqRNuq8wN9IQPZYkNV1N07
BtfqEzOMPImsxJmBxWIzjqA/iS/5rgqTm4Jf2wHOo1QPvmU1IbvTUr+kbQURQGVQ
5fgqy6zmMrY5MJmeh6PPtapW2M7GF1LlE5vy8bHxhJDt4r1LNDvWiCSL14mdxG/u
OyADpZIerWP4PdJNXZ6Vis1CUF03KmjEIzHreNLLEdzXIKU1IS6TSr8cQLQ/zYuB
LfVxJlzWngFcVG8nMYBX31dnMBRXcOnDGFwYC/3eEcxzEYwJDEJ2E1NeiLtPZV5D
UMM0weyKg1yTu7ZjYYtZVE2aL/bdh32TXdtlrr8zrXbky5lu3XwbeYA+79pWbcMn
MGUqRU/igmduPTFRxRi30fxEMw1OAGu/ZEbbupGmGyNM9hu3Tx7XZi3pBpLtJh5L
ES+3+/gMvq0Esn+WYgSELPyt5MdY0F6drbBfac/e3g+y70XY2wdaAev47qK8LPkI
nzVTVIL4dIZ0Tuv1DBNMC/MXgNL9n6xJOhqTOiJzSTBcN0M0HwYROqxcqqLDbCXd
uLLy6IAKAPZVilTR9b3veYMWaOyw2TN5FQiSqipwPcX9Bk/f4NHrxrQ20uYnSdjU
IlQ2XFmrkoy4d30zRWlKAQWWRh3C6o3gW9P+DkaKcitnDyKmz6juQ5G0r4UQqVPX
iu3Mgwkmac+dPZhJLNfWQJmVab8X24iacQO8SuRx0//izySvU6cnCmNDx+Ut/PNv
zV00oh2hRhma0mYjb52pV0H9IHa3SgA7vxt4HZtbGS16wf2NOHnr5TwQec1RVnK0
jmytHdSIQz/Op0JMOk28PRL0PBUz2q5Hau3PIv0e5cP4eENyFXLfgh2ytRr4kcZi
aovxJVmPg3L1UDcrFnv2kp3TAjMEQnQyCzjPhCCQ+q1g/KbyfcaSwxXj3lRL3PTT
Ut2uIQB1NjCYXmDWFZKCPHJj2XgNDQu8PwK5yRW24YLX9f8JvBtVuXbL7sCpjW2e
rhBfG3UWG5A0r+ZUR8uheozVQeiemgjtmxr3Dq8L0RZybRYiI0QdLEiplj32js6c
/ZsCEdVZpBLn364TM6VQcBPD45eJpM4+ClH71YtIgKRV/Icpj4gJnilL+q2PWU30
e78YEAqKT6RJdaVfzkxBR+hVnho3r/qEZslB7BhV7vQF8mXJF0HFZ2P2SZWKAjN3
PL+4u4jWYAHsGwLLNr7/+o+vvdr66efn/1r7jgFTT4NTlALxbqw/jbTf8I3KPXDb
uxS2EmaVunbcTIxcRKEO3TrCTfVbLHLobSZuS+3cgt+cqtMUk1AfdM+DXfA23OtV
shsXav4fQZ+FT5R7A/JxXLowdpJEp3jTZYoNFo9Ik6WokorGcAB/20ykFOOyYLvB
Q+TDRT68b92XxdRU1ZbjiDqWvlQP/Bf1DZyc0y5Iqx+V1BUqvyCH87dQOz+7vPAJ
G2l3bSDCQZIXEFGW/54EmRHADczQ1byhhGlfqkNK69qsw3x+KkEZ4z7P88rB1bDQ
SnuCbTQNVENqRi/ozr2aWVVFwijJlzbDPRUT5js8R/sdU9mZO+Ts/jaDJ2AZB4M1
w0SQZWj5Vc61cGkZ788l9FMPaZ+RJpLidksVT0hSd55nFzzqv4Kw+Cw/VfQoQF/S
6DzdcaU28IxpQoeoFljrrS3NTdep2hiGSeDjZ6yVtxpLDFUCh7FkM6VlxZaS3Q5q
uKRkREXjSjCEd1QvyQCoy1mQAgUjwPhSO+EiN2dT2Ov7ZD4IFKjeHsCR7jkjCxSZ
OIf4KMFh2xvM37OdHHICj36X8AG755sYGSx2tbzqvNWyn2X9NYg6iuXJb6B7UVfN
3BMs68NXcE2cq9MdmdnFh2cGr5tcxauYPUHKBw16Y17Dp54Flp84nxFOw0YJs4mu
39lKCI8I8ZrD32HW3UKK/3fJg8F1+ZzIr29SHHFrWmYe9Nr+2Ri9upWmb6TC+fdk
bCMVHS823uAqjWrd1BonStQ2Aqg2lOLh7ti4IKnhuERrcNX7NFrjtcUdqFoxJylb
mhsIAe7Ew1Ul/UJa5tzLtYHjNwJ0FOSkObPdpmLn4fxymi9Ip5rIzV7xzK3agMRE
ruWj5wWhuYdwgp9Hye5Z+uk0KvHUcZQ7xjSTLt17GDTwL+PzIlx+lV/wLUfIUvuR
VJP2UUGkfaVfK0fl4bvC+rusBsR1hoD94GyBkK8FP+9MytjV0lrEtxqKEVuNZnq8
aq/lh7gV5GufLnyBIBVi2ERpkBX5cSWvUdhFjIm9QTzAyNp1IJHwktTMkQZsCERn
sf5+NmXHMP0BRino7YmwWC1nFVJIcVg1g/KvbV1GVU6Fa1rSzDnx0qY60zBGqRlA
ocruN+fMA5TPJv8PgHNur9hVNlXAx+f5CO95SiNVJFZiBEq49vN/4+6eggC90bQl
E2BDKwoWT9ABeGVIWGcrXp5e4zcmY5hkV0AbAQjAe3qbP61BPSEUhbKxWX+9od0W
Kg2+F6kOXKTeKBCQeYCPwyjXBKaknTWrncFTQg+j69pKa6g2rESvLB54Z1ONHzMo
DPGgzLrt1eR3IDrGfDHso8ROLa4/vTDJp74X/ArmCRRWb1766WkP9sGHyx/ISCTU
elQ+JJOaHfgkVRWiW86eF8RVIpzPX+43XS2qnGWKXf7+JxTW7cnlvqQ2KACikefQ
CMYVkodNTM2lfgejdilFqbVcunrEqQ3Bn1lDb5w8OgYABoasQZ4+zCk8DBOQbfZR
jn+FxdC37BbflvPmURLfdzcb5bppJ9Sj5Z5ZYPmAUUuHNrhz9oJZLqIvtlm6nQQx
DpooDYg3hH2nnjvG8P8CrdfcwgXCJRRPH0/FkCbw6g0i6fQk9DQXJnKOmxa4oaq4
tWO9Oc/wLZzm+9vyJoxtwsUHzWQ1miDhbk7XSfcYPSXAHz6R3nK8PZ2+dJ8DDS8d
pY5e/tjNiRypIXLqQMLaYR456o6pqo6DXibTwKqQjMJrJB5rLFfJMsL3vHEJhAcH
abUFwdkQ1dNCL2paZa6Rs+2OiJYoHSCg/7QG5crdDgdHpK3/hNtgtwkE1UfWAZ7j
dRgwwWr17htmylNnmnMjVmUVUmZ4fOc04FpabpY9wA9FjiG3E8wuK7tRsyhUyuQJ
2hIGKxJAF810s3n5YklTFPlab+nbj4ZurlcICSzHCkrlYTFlMUeYcCAwsfbCZVTg
T7kMrj2XrE+99OzPplqVD7Vj/cQDzakGukoX35XaLZT26RF+u6JKiwVYiLykA+mO
cb5ZhbZAVHSSHa2eWWlpHtAy3UxAR+l7socdBhj0P2oT9/Czm4+JLI9EEijqYyAF
KSczGUTOUIIP3xE5Sn2QiGv1IbS+idLxtJeeK6g1ROgpL5PX++XpfG+dkT0te8H0
sxIjiVLD0xYtyYXlyLPSin3yc038Q5qImHCnAkNFxNTUO99jhn3mc27CVz0bjI94
egSFm1lck+MgAJPHh40FblK0AO0F3yhTilpooNXQTlayUlyiK3nSUoBEbifiZ9UB
F1rtZAIcvrdjpELkw5KocnfsSucBri7tTqYOXunjkco75AkyGruyMWxVKSNekTCg
1d7iO0nX0JPtF5pHL/Mx3Cla5Wl/B2PhqaPSiUHHDf8ySkKVgeVdmOOhs+cMqYgG
LGI7yvKiEOE2XZm3f8BeKePHW5SuMDduItF8wTtwmEJ3NgdAN2kCWeEEzA+pxg2f
QfGirVbijVn/QmaBNKEyLi+n3N1eDWM/dec+UoxeEBHIBKhBBe1QmqtkpzEBsmX/
VcI4oniNrOyM4Y9wY56h6IwYNq8amJG7oUUgwLYpPjy/0pPPmut5U4tYVCsussj1
vuOPKR+s96FW9RELd4vVZ+vuYOS8fZRf64xw5LmSz5U0svc52gdqcOmWouISLIpl
Ofj3i/L3DVTMg5X/y0MTl2j6RERCDzH5CjqkZoJnSpvqnPPvwxsbOfVDv6dxG3Yu
1YPLB25d+FJaRx/mG8lmoA59UqWwxUHfVPZUxQlu22BECKE1u2RpqXfeFr5+6j2k
+h/q5PYw2R+XjvbNjvRC8w2vzSbv9Y7rn92HE6SPe1mu0vYoEPe8ZfY/5bnsLSEx
/QSoVsrKAZo/Mz0ZKSyHnfYxwb94pA/Oc7veOTZ4hKdl3D7VJwBGmJz5cZPbubDG
W2i9lQGobqsq/oej/dkwj5bLumzbEpvPRihnfS5XLJJ4JWnr6XZVuXFXqtlJ2OGR
o9jEMFATrxBQcWDrlgzvxsBNcEsQ+aceuEm8imG6OPNd4u/Xq/sh5DUK1MtVhmly
xdaRH5TI/I9M2xOE1V84GoqrzJnzyySxxlBUZDTucWzCP/XayTCmAW/U3TljP3WE
ICQ5/wybnDSv2ZSLQCmFHeCfdnSMDhcJCnifFn7Nc6Yg61wUV9DdVGQG9JbrdssY
3HuiurGq4dLqv/7oEzEM0SQihqwwPixvrgbvy8vvHIKccFgD9l/buRpy4uT5HOTG
r2NVvIZjmliqh5E+rubV32pMdi5SelYmy2rYd1zTUJoa0Z1IMO1AuuM/ZUFCp41g
6pEnxh6VqvQy9Wj0yABchC2QWl4o4wtOyMU8jz9ufctEC1HNzCrwJwRLL8zlBtrc
0JoPElDKVoRN2/W6ruT1THELiss9hdN6vFrtiHXRfxggs3YyqEZcdEW5m8Uux4oh
kQ0aCpEPiJ4EFbiB2Eywh21h0sAFdiOMId30zjrIxZ2vwgZRjJdce4CTmh3IhCyu
I/OBLsizXT0tG5M84ojFmEz9SAVGMvGCLRC239V8pxOGSMfhwa2vuRtRnwy5cYEf
Mhcb6h550GXevA+SbI4v54Piq4RnJ/viAKPdbTX/E/BUOvyRzJuUO8Sm46annPpU
zedBUtxPQzHHbMWHlabxhlEnJhNwlxuclYkScKWKrTEVI/vPmK6hkqz4fEKlwROP
o+IjYBwLebOgaQTfORz+OE0qO3quO/c0+LksjjSzAkNVN8HjY/1A8/9R1RQtYe4p
FxIZZ+oqS0ioPMz6167lCE2py575XZU091uo6TJpAICzJC2qoU28gA+RG2usqjs+
uTQg8fPgRx33lrtp0NK+vhvi3xmGOG6+pnLkkjc/O5BuGDklqbkYOXWH06sWfZlT
FK+gQMX0px4xcUyctl5mNKMZNx/nOfYdl7j77M3Mfk+DaMruDtcqG5jmiB1Fqs8h
0W46/j+VD/1BXgv63wlTy42USiehLhKIZBztc5Rasyqvx0f9Ea0y7fKFoc02zrio
EAzJBIAvE7G9pJAuzXj7TEiKAV0Xy7Be3Rs46PbmLrFNXhoaKWOmPpAWzdaFekR8
ckYRYAXTtz3zIZlB4ZZwoPiA645FZ0tvWZ7wfQhRjahnn1QxNdrHH3huOMejKgRL
Gm//vtK3ATjfR37VA3ygWf9XtoAjzJoG1OkuqvR0M5O7pkEhLqAAyOdU9da3uV1b
0EEDT7A7P3s8xHWgE2EbODNKtljjjuw/Ib6AUYj2cZgsIaicaVxzBI7ClwCPCwDo
2emSP9qj3kkMjoOZ+oRB8qP6ouaLcAHoauzx/hzD/PtLq7E0bFXBGx95/I07ynUu
QAcPZ0CFGjrm2LtMz5hetW9SaLlIHm4aCSxVPwOMA1LNvEaGVFC3qa3p2654ulBC
zCNUwBP+fghIo/5u5vxEjwMFQ3kB0tjmERX0grvk7ViIFsmcOhxzhDT763Bg8l2R
3Yc/aYXl3zHUT+FCqsLAoMwY0YXPoO5NjQS8LC3TRAEcOSAISrjSO6F+R/gh5McK
da/nP59zZTBLfhixT8fKGKpeOovyIyae3+zyx6j2bpF8meYsZVIJAwbzbTNfq6x5
MPSswTQCyjfTEhN5G2UwR6KLXhhrdBljtOiz+Yvi99ZmlJuq3RTYbxVj82RRsrNp
t06GEkAVB1cOam96O9P1EmkemFP5L7Cw0tL+0QnnxX7EvB/ZGdMCfpGF8GlkSxCT
rluUzIervHY4y7O3A2YJPVj9CRDUh1oeXGnaLmAooP9HFtFnxYFJYuDzUQJsW6lO
Cm/6bn0wGJGG8wpdfgPIlA+NOmjHmvZFaINUeE8qifwmstYVZEojqSbMpU2gQh6W
LyBrfKGlcksPAml+XTUpESHdOHi9RrnuqLBTJHu/kpou0pAlGzoTjuuk9mWRNuS3
/GdGUn1RRQWYR2Sp5o3vkRMBpr5eDirNXv4G43nHVFCznQYdZkbD/HWPLh7Phzqv
9rwKeXju/c9NHqvG4OusuULw5McUMYaReBIGKAV8aS77yaiJyIqbb+fvvXW+cu6b
gHagvfGMAA081Pac4yZiG1woPFjVQrsTA0kLidKbPZUeSm5lo14RmijOjnHoxIby
gutSMrxdWc43PhQ2CInQPdHpmo4KuCMRsIlP4ltIZSZIf3equ8IPiXo/KFUBR0kS
AZ+RnwLr/4OjKehb7ZU3/bRLn47pv8jRQJ5CCIYJZ6sVEuxNpOpiFfLMudhAlmbk
WJjOE+VzEc4bHCv4W6ZEghzES2EPQ9AB/NxNLvEk0LIV8mVHydjr4DXlRXU9Vcjx
1taUp1RkfO32f78fBHaPZzIb5LaO/+YvlvdOmg1l+KmsBp84kLbm3IH4wtF3bnke
uHzuSPqoXqnhAzd8uP1kcsYQDX8UmgZi/2UInqN7G+vUOxUMCMCshi9HvXZ/do0a
UHikknwqw8Q3ryGIieD8D0uYbJF9C9xYKt+B2/iJTnPTARpWEpwaOqwHnUB8FapG
GmzS4u5135yrhlEeiEi2dCunQLPrl7PszO2lZlfmgv+4O5H2RYDhBkU4kQS3YcZm
5fTIF/Coz2IDPrjfEjVvDc2/CoBT7fx+4donxKrcRBLiWv2bh4n/ZlVG4augbt13
lkKd9KerHcI0xnP9zTNJdOAJPQDG06yls2G5BOkYJ0oiIYTpjrUgF8H+7gD7TcU/
HmkeXqxGn9ulC/HaTNCDUqiFLlvnhq6vYLGXXHyZaK7WqL1ZzmqSIaqmHwlcA+6/
IJyTyHooXI/5J9Cv8Mj6KdbDM38AGH6LY31W4aWoI036YIYcoYC3NYqXP64HwRs2
bk8ijBf/rDTistSEb65vRTr2+1I/wUGp2Cvk4yh7RAXx1e4nBMMcBrsNjkQhB5lS
sfXOMN7PbIs5u/814dE3UckRA6ZUEL8nnYUxWby9B8Wj4MBmNZCVJb11HQKgvBBs
ehRF0FzWJ3T/WKSXxuIZgXs1eyWOahkBHqMhBKQppAZT3o8b5BuU/a03vzF2tuvH
3Dbwn6iR+D3ewXGK2WEaMEessdMkU89F+GwpkF9y5JK401pl90YH4lVEZDD1CesU
bkZl20ysc64pYW4lskL2rwHITDSa/8uFHdjTUY6ArxWGC7kH410iYIcyWPayoJ49
mxpkHZ2zGynBuUyYfPI24FsH8C/q/KKqu+6+M8/1IH/SWgsY2U8HNnrRpHkzFcvD
3h04Yi/+8h1Un/2DNJ12lX9q3GewoAcKMxU9Gn4nCK0tp5gQrTA3G6f1OVTuh9zv
0LizdJ7WPI4dl5HjIWZ2JJ8Yi7r2+DrYK66jcMklH643fPkrI4d+JEuLLK2M+sgl
/1YrpcDk4FAgqlT0jjz2I4GLPVlVtxF2X25bBXc1b+nV9ao8C6HeSdpQ7m3ZCtT4
jio0lKh4JfVR3dMg8gv36jMH3QGsGUfmnyA7d08pzn5Q3ye+v8qJ5/pKT1uUjikd
MVRKPH6KJmQaz6PmCMl8WoUhP17bEj8p36KBcGZ/r2JBczw16yeAJzyCtw00tfuo
ycM/s0rDsCnAK3xgJmeEcu3XenA7sRmk8sKORfvcMRaUmklOtmMfEUjkm5R4/rIq
twOFAuvxHjaB8SQnGFe21VtBlCxT3R1Ir2B5UfBZi6bThBmHgnf91Hl2seDKOCEV
JrhTGeHzJnNHBWZran96UG8t1o51TSYVtfgpSPRfnN8SwtY3V3A/v+XUl2WE/Nom
PhfrTZVTa8FJ2da7F6pMD3amYwajhhG3Nqiy2ufREoV3tXdJtsplKqU5bCcZ5+6E
ZlfZLrG6PDPL3ULQHsIz+OocAMRoa3ttDPIc0iE3RQk/FG0Jdx/d+lA5b1ox0j0I
CZ8tQjb6+DMgn0wZ+JGF2bk1S5WC2EVzOzLRjdAXpprQ2GCK2cIsTSVdC38hJRo1
IP8Cl5fI42ps21rYPZ4dVbarq63fXv2okbCqAGCUeNhU4zbuUSMVV9oM38WPibhy
NY3vQItG6gMSxMyhVqorSgfW2sJjO3p1lytO2T5m5I3pGoXJ0oBIqBBNNnBsJY4K
h12cV9znIGLOJ2DuqazmucLpNV2D5gP1oc2lVpuoYO6qh3IojpWtqaygKbAoItkx
J39bM9kAAQVeGkSdnvvFpgNzG4hCYCONtfTtQvpvtqpMPGg0BdtLJIHzvk5oF1p0
WqNANWn2BqB22awzlnKwzy9JDz/Ik15TqiPatR05QcyYJDcY+4sD9jQsorysAt27
WliUJwen+r4/j7Kv9YOj+l4M3bzfSzamQdH7EY7ik+cOygY+pQRJWfVKXX7WbWxA
d/RkF2n1QpOWxgbgleabnf+17Nc2Jqi7kyJjB/qc7WmM2ISfcSVezk9O61nTCS2/
Mhpl2FOvXXtZebElO3ui8wkop054ECSx4oINUvkFfMx1RVn/6J6TBIaLQRGw3nHn
N2Xar3FKUygO2MePVnvQyMfVkr1kxAd7eRr8LxO+1M7rUhp7Am+wm78MI4I+rXxy
Q+zpevG9/BR42XGwah37NEuVzB+gvCwoj7XeLsBnCq8s4rczdh8Sg2/NU/RrASpP
/58AnWtziKXp2EiqsVu7HKIqsa/LeN0vw/j/458jNw7GNVzcevhWb964//QnLTuz
T2sjj5/mhJANYiF/lI4hSofdsXiou3nM/F+fCmTrJjFmmjMNqs9OC71m1BStkZ5d
Jks0JQ/H+dsWRzTN54e9TeGn2Zb4loiYgrMiN5UEUKTeuxmUdVl7xdQp7uIgsp4/
rd7CfX0iaZAnrsnphe0FzCfb9+KDFo8FjvTlCTHxlAy3a3gyeBUvcIibgQXMbLX/
2rcBWZ5wleOF7WP9ydvkSM6GQah7C7BR2WAnt04YYOIEOXHw5RTymWqm7ClW/G3N
KxF3gzK5XrWYJXgyjSPjLle1i76W/MEWA0hBU0mUazS+5S1JvG85RMgr2VKtelvy
x+OfvNOL2bdFd7KBbTExnoF+BgjSU2wFaUoThiV3RBLCBZswm/l/FX3lsjMqDiGt
lqDRpse+Lcr8fhcWQZxBMNSVchXBzFsCKE3rN1ip2bT8Q1GJ7/H8sgCsRADiEdkk
/O/wsXyzA23FOyan9b6scLxRvZIswKsTs0kT7lmIO/fAkMhSMK+a3kbsaJ+maACP
d8angG4pzDrjfAodM5JoT0H2HjnhqXjR1xpl7daS6/uSTSB9Pj6NzlsvPX5n1Pph
OuQzbGInxBB3nK+zEA1lpyQXPpegFJhcFECTOm7+N1zfLRieQ4Q3qf2dNwu7lVOE
7/NIMHGOGV+gY/3AzAQvo4XwoUnHGUO7in9WrPNjBhvD5DK/Ub3uepOGggfXCpQj
ilMbtXXDqlhH2ePpoEcCLbgx3tRMg1Skff9XmLPY/OEjgsYaTHyBV9589Y8pMnRK
6Y/5t/sCqJa95IA8md+tZOe8THZJQ2eZyrFbughnRC5C+tJZOcdK1MK/0Eh4E5DM
2WaokwfV9b6Zw7os8sr2svjaDTy+Zlql9yAVEEtoTdJaG6TajCK1enLXSCgVXXzv
xXEQOWrwYJCoHK11DmO5iZ7Q4Obfr6zRAOMSVxBDDu6cApHrh0YnnZB+kaEzWNTL
nWa5PdE+MLXbe145h4pu7shRRLLospADGq2Fkq79KE5k+vXOKFt+4PpiDP9PAkKI
xfPN5xnVHG8kToCKmIol5aent4b5h/GiwnAYoL1D3VDVMTJFCty340f1WCpXzoPm
R3XdDvF2KsUwTtfh7/KdWxc13XINGhlZqxBCtrgZMTz1Kr/qw/AeQjaLIgQCR5J2
go2Le8S9oYdyiUq0S9On6PTFM+M3ao8QjLThMomLTpyco7bSWHsrS3IqUz/UpeCn
ip4VX6IMMmjJxG6ZxhZSb7l5I5I45+e3UTobeY3EmvuYK5acF7SuidL57sU8pr9T
0dmViZP8k4xDfHIX3h3y6vv20Z1gRszou6zl7mQFFXceyBqD7OFEFdy0voAo1Lo0
8MpdpDZGvINgzersgx2n4sAeP3UMAg8iHOydLtdP9h3ZVGpYI170O2tubP18tRwh
p7bC58Tm69qlgKAATzu2EXtSPa8C+hleRcjUZekQ1Zap1tnrjMXk2anowJCgRbvJ
FG2Z/niVUcd+g9asA9xaJAJt7cAFtnL35X9qG9NZHytIgm+u0PMEij3KBbhLpe7A
XfvSY1N2YEXOPzrMkz15/xzVCxE0l/0hXy+PMpY25V1OPhcOcYWweMhRayB65ntW
Ec2eLzgGbZjuuK8FMWr5KMOXBv56yowaSAm4DkoHW0G1+hKxcBumDA9QUCoD6ILZ
olp3HmoxKrR2tWG+su337PzVRH5NcZpU9DSqZcZRC8saNdOBF//+ajVE9p82aZM3
mE1hDzYemJrNlC+x9Zbp/daBLJfM3zXZKwoCnFGh3dLKH+5FEOEpLFoH6UqUiUlE
F7C9KKC3u3tJWT50scBrLRoXOnH+0sUZw5PkkLdbdt/NXKXYovkDIgHEx6/FYcfI
gGk5bkuqky1wM1WI6sZIiAAWUUBNQ0nx8cTx3t/w3Q0FKTIJVf/KnHrB2OeCkDmb
wbzEDWTOX5HXAouBJ8hCjpi4O+xwOkkJl1AMbuyw16GYFsszsad8ZAoWk+DCwQa1
Y/EwcuUD0kKO1XEfmd5a3Pq/k4hIUS+jnyiKZ7bgAOdYWoxrqeOUg52en16XEqfQ
4zUqi2+PrgqQWGTQqV318UPxj+nPaG/t9hjtw1bph0ICIky1g8hvwUgL24m51zGv
0ALOjz6ge0Z6F07m3QtEGxyOv2CuB12j6x+aCHTsUxb5h2QEXy3JQn3vVSIS9bnu
HocIRepaPJPekqQPReza6zybkPfsO+/5vODvV+SXJQNzMKN2nKB2P2NVx9WNRQ08
JhnaxW6g4ioYLDqbxpqvxjvj6zGtZLuDoUiw69iOWkT2oG5fQDBlX/hb0+lEApZ5
TUa/FVgAQRtOol4Z6h6cka5z3uNadffUBozPU7dzVK0M2AlHQgEgPSLAZo0mnfNo
9ogEquzoePv0xpSNhyUA/uRQ7r0biR5ZR4jD2Cxo4jwf9XtEMG4OeWCAYSWH1ZZN
7v1vSLI/44+Bd5LiI+KXLffr2wDkHPhkBY2g6RC9P/+MHsPgR6XlExYb9jA0DYBk
VKzgAHEzWxX2333D1s0eoy46jNg9wKHqY3SNM8kknE0gwQwrDhy5Tws9wFPJcojH
5lbAkeFqpqOoMEa4+tYCgATZB+lODYtL0+LvEfmnSknGNFeH7YWLTLUyQr0iR1Jc
dgPU+Z7kiTie8QfW7BnjpCaKx1Og8RTNu0EJ/nTwTop65mTiaPbXFCdB75B5gpIg
AOwUd/uNN9SdojKGmvk7o4eKjc5vJs4cm5a/eQb3EG/aurOTAV9gvqI5/EXE6Tzi
eI6OF2Vi9m8aVytSx9kVXytq2O1JXPxOYtK3GtVRnRKMRUCuC3UoeFNXvE0xDmNT
n8V47B7VWftZSY2OFfd4wS182JkgNiTboX+INIHl5SZixhInlhjkjbkshSrHBwq6
cSWbiRtvo085Ls/80lfUopgfTr0/gq/Kh6cWF2qqkeFS9LJfSmHBlUJzmlj/gioz
ldWjazJlMRv0HPFzwM75/T3Ro4uQHnc8o7zLqATzdfr665cNmD4iUTZE/Hw2PgR5
OmJC9dK5ijsDZp5IBBDgQlQqx9dvVk9jcZecLSdJoxx/iS9zRoo2J/tliV0c0+LY
q7M1xldTICV22OtIuF18pL/62HnjIDJDdjLNdn23D4TL499IQMMelNseV3LTvYLG
anj4YvB6eDuBWPE7xVAmGWLqSlBxtQvNLHgK8vYMkxEtf2EONKN/dQEwnkUnROJ4
KqoAjeYad3WYWOLAUU0oH6lskAM6dWDKsAoSbUFKZVMNRQiy73nb6yikeSPJWRpb
brIM83bDApTrIY2PL6iH00G0Yu6D74dOPGNLFTJGkdAB2vCNekH4qNHgf1L3X7o7
r8q3cVBFtoHgOVZ4HtL1bbpvP7KpbemKiAjKfrJ96hb5+FUnrSMATI4KIS4Etr59
0kmiaqe1B4fawyGbRncDrsRZ4xD3IZBV/rehpLdTQWvLlT7pXVXU1x15/qSZfOBR
hYgymV+qGN8acOWYB1b3Kac0CB7yQ5KrnzHOYaNLSNUKImIFxmoQCPUMHnLQE0Hs
Ne+gsdHlFPEk6BGvpPpBlcuI2AODkPvGDdAz2kqWhM6kRi5BjQBoHhoSh5gPXxSS
RYiBQZhbuNt1O3+eFy2Yo15ieDptQPL8QOmZVMaOGvsDeFqFxY/+56dVjkSvgXCK
KXUOwack7xDAvHXpFm4gzTfESVca0oxL+wk+pzW0IpDVZbxbcsBPSwx/GfxZIUcv
QgLTXvOkGDXPRoJ7vQPGA3ehSa3vYhESUictSXJtTfWqVvCSbhaYM6U8Ht0ev15p
manm/X17Aji4oAmoEO2STFbr6dNwn7iH8Cd2CSHZujXr/cr2FQfNjmTaY0hzbodR
HPGtLz5DPAx/qjyb2L3PDbLbCQlG+LL6Vixk2vjmNFI8MvtUu0BiWW7/OJAEq1nq
J1t6p7XyFDG+cBF3MVVIBxtaiRv9RMloKWoWSkGzveUGYdAs3hHQIi+/u49aXdfQ
UDUQvoPgigBZfvyY7LueZKo3IBQ6p7jyeOVTmS4vELLCnA9/Jh/d+QYqq+kBSASG
3KVgA6hIlD0imwAr7BNf0D61oavFGV7Tcm18q0pfsw5b4TRo7lVaDUbAgovSSL3c
edAsOvfJAy4vDDpNAvxO8UjyMgf/kXF0aUhxVlnKTrRGMHRN7u3SxJpeL9uqjsRt
10gIQb+GllgX6rbv3eqa8kZpc/vTTBWrI/LGEvG13hKxJBrit40HD0xqDhNLQfcJ
xEifAiz5c3xNuYvMhPffARgQWbDBdTw7C6gyX74gj5d+Ih+fd7xVf3G/xj4oaM9F
LN5H93b8Vab347RHhQDonA4wZwjPLeSMN5ZIAo7Cx/BJygY+balzb/pB8yGmCFNT
tbrcdkFl+BTJETyGw1Rtq9+C5DBMWqEnHqT/yX7x0g84q6k9UekuP9DkEl+/NFPP
ZZ0QmXg6HoXarU1Yyd8lv7NQC1gkmdsWlYi+NbUSvMqDL2J8zUNANx16vmrfznMk
JrjXfA16xfdI4Yq2kb+0CjZg/IlRCdqgk3WHM4ZvkMDGTlQD8Cn0Lzn1E1IpcLFu
N3GEs1zYP/BpJIrgohOz/dBydPUriazsw/XUnXAG6lkWag5Afdaft/gVon2J1ZCS
mvxPbkX5r+SO92kmDIypptonVHhA8pSim6p3Q86mEGyU1pSiYdEUtnqXsK0k1P2A
xM6tUGPEFZKVFdHf/XvcivjV6gDFumkShk+uQckSvApiwmvhXLh7MytzOeMVf51M
pC/iKvraDdNqcIljx+YhM87unPRyJIKBg13NGWcY7p2WDV5lKZElX3YsVzOKM+V4
O8pRvn6GbrPJUBQxe1q517SPjkt6rr8mbL8MvILEAvSCBksqPtiPIB8yetd5Uw3b
l7ZTik4Oln4wAir20iThyssgkCCaS6QMIBVChVMWWoCQdDeBnxxlY1yuv57rV2V9
iOtr0sMlKBS4kIglOcV+Ot4MD31LZR84sdKZyJMMuG9Ig7L2CvtIaQS6GXmHuikk
1JUM5Wcat4o6lu9J8q4nlKxiuY6rqVtARPZEEOCQsP/naYfDKwx7wz0/SJuoxZj0
/Fi91T5pSPT1AkgmoznMqx7et+PbR0sVcSzpFlM1JjoDO/FRCzYW61NkFj2nezGK
nuxP+M7WMGs0jsyDIhKztt4AW+pL/dqPAWEZt9M9M72qAZWm5VYfAaWy1d5rVYlk
8OICq6oRge5difH7b6GztY8UnTxCtZdhs0rOHe/tp9CzjeZpNHzd+SUWgmLDF9Pz
6FmMKHf+piw4J2o2cIprHHgJk35mdabK8ZbjQEBHe23B65f2bS6DiMBS+8RK3lzT
mv3zqpNCPoOK6dWn+Z/z4KPEIOnhrWiAyXIdBUrKL81n6GhKvaGhw4y6XZ/GM3wh
e1T3gUkO3eUtFcrmIAb8Bi1OViLifXcLMDmOD7efsBeWyCFKXoFsh8Vluu17LQWY
eNEuQtu7h8s6QJOM1vXq/uGX+oGHSDhPldGg181EB0lZ42wLyT9rXZozpcpeUxbc
/KlJFs/rUMPzLZxeHVNbX3GFVVniqy3V6FxN2B0C71ZdsnSSWOhmrx+d5fDiGhpo
9DALxpGiP0HndifpnO25LBYNFQ0GSIJ3zSSjJMkrzTcVdjLI3gwbb8R3DWsq+npC
d4iDE5kacH0QVBoh3H+Gsf45p+/hPsjbUOVL53vCfQN+q3EXWfAbyuSiU0bXSnBV
jHFdKhIwB5gOhV2+MnNkJ4K8/lybjF88QlUoL0Oh7beTH1glmcC656OYl7qNcvTY
lg5nsK/MvLWzs9HWph0pfQGE4P5evCxJae7U8vlLJpmpixVmwFwClbKPNC8xU2ot
vwIlvsmHTsTVfT1CNBocU4b4LE3OljS03KN3rK1pJsMOjNWwDycz6XRGCFranphE
ocXxxmVJwMJ9DOAfrSvEh44NvM8kejghWNXpUFCR2w6ImqenbfGo9KqnJiFDdMUi
o++NO2TbMFaHlbPuEt+AWdLqS0KRAlDHRK88zszwPRhKR5XGSKOr2FDSCWsiE0ab
5id8NAakiAmuWDXUQfnYYU9dfr7SqrVeR704/PYdEstP4RVgNnFjgTquwmIhnfO9
gkhAcF1+Bxct5hAWAhxPZAHm1vgWlRR/oUQO3NUiexAPX8A68uNAZlAfMyxNS+Kg
aomNSwlGpLlkhP/X0ST3AlFgkxe0AdtsP33jeNGotG0FwEt1uX4D78CVGkh3nC9L
mhBvUAE5z/NGvStsDqfA0Y4/6lmvtEyKVrMXtz6iE5cQ8yqoQJKnyvO4raM2YBhu
w8mG5EF2fJ9c/PbIpBNW5NWoSPMTK632GhL9qTB5uRO80l61lfHUa1EDrf54e5Zo
WKPf3p7VOVUXE97GjJatO9YVjPA+PuEB/6ZIdTj9KBMmUclYiTOUFaqh0UzDrAF8
l57NPasXtD6TVIzf/pwdZTflbJ6AaH7CwYo2zloF2+s9Yv4EAUHNrqi2v+MJrz/2
WXf5FKJQwvLcIXMpKbu4FvmuKOAjwO8TyECcRR7WHvrwN4ZBXg307mkU4cDeEl9r
en/5nk5QX8x2K44K59hi513WiblFydgUXb6MsW3gg6wyrh8JmVjBBClZ1AeCqHTp
oVOWgZbAuFouxg+P6cnNe/BD2kT456WJ8xWYPVVFCiTSFugnxq+itEP/5fYQCF08
bM+7y8z+GrywwzOrBGvBZ1d4SfhrWEyzw6zVsIOp4J444yMZQF7tJf2NkAW9y3Az
RMs0K4YaDUzRr5Xno7LzyOAqzYG3AUe5ZrSvwYsGtZYyiwsLgKvayYAXltbui35U
ynRL3UoCYhkYthe54Uy2KF5dyy05dATJVYRUXJ8hkmlUQwEqpTfav/7eww3Madsw
WLMkqgHezAIjjiUDo+iQJgjLXldpX+WWYiGslde2tUAGi6aj8HpNmLyOkxJ6r+9P
Y57Bzgqwny+8XSEgLmxPSKErddhT4D2KPkFsPAvfpleACBbYzu7bnRGht757vXfF
RaZWWQgBBOLvId8hLQOJCeeTHOsbYOlPDc/l8FgSLThwHyEdrFhIor/KgCoWaVIy
uSnvbLEhLdwKn15kX0rpgjmU3obgFgvOrRGEoQ7J7hbL/KTFLZtcbB5AyKaqG4qP
a00+dAcdsfnakbJkoq/zLxnKynjRvKir1XOtOp2faR72Hhd+HHQPseFpU35/pUOi
xeNXGvgyWvxs+Ry61Pcfnsw+GUWnBIW+sIlfLYYawK0k70wzV/DI/VHcTcxy4cli
MK08mdSrzrelkz+6vEF9Ncbr5GNg+e0zbCi2KCN6Ea7M6JvFAXkJ0sEMJLclR9l7
TrmUv1v7q2xZGhFYRqkpDPspagA0pUh4HK11zJ6hD813F1rroXpEAFD25o9nmCcz
pN06TKHfq0X4/aO5gW5KonigCC2dqSPM/S92vU+dA8QXNox2MbLE7W7PLzz3K3zp
6nyJmijsBXsjMM2QqJasqIJSIWzfNhAK8W/J1AMD4x8jA4x00fLmfDIdJa6Oe7Xy
8vPWWC5DrLL8c7PQ405lD3TnBgAlaudHbVDC77iPf3wemunGYClK/f3YH1H3xlo1
D0TfrvRg1F+euUY1HRyvzC1xakjZ+Pjj15URBZIqYjkPOUpsY8m7B8wwOg0cbkvn
Gzk9NzXo4wWzjtGXih6HXyvnsI4WqlQLCm7ZOGgURvttz22Yksq2iIRqWRcQuXpx
vKey2MGEnig6hZJ6hEgG0NsAmQMSCtQhXFk6MDGiOFt0JNozQUuP94DsZ36mhULe
18qh3t/n7MWQEMmPjLsm1D0T3ccl24dANFEHxJE6Tq7/3hO7MWahixvBI/MoaWeO
DG9e0IqsYz85/gjBwBdHcQOvtO6bZk3bhssj5FJjoSB2wU91K00UCXKEnNZMw+lF
+0UMWmirpecwegTrigRjYB9sk5UMQ8gkjIxAp9vsVYdaLtRI8tCLXlzvgMRfUJLt
eUWSbZ/Me8Um/GGI/q90GPAm0Yx+WcPrbyckyn6Y4vqH4jkrPsrFgwAXhky3YwS+
5NZ1OOVXfUHqFdAqSTbMGN8oDBuPfUbZOqxLWq9OlDCSN8EjzW5JEPmW+q7gnHib
mTy9SX5VIdqYfTPUIJp2cnfYk/JOfP5/SfcflZxCqtwAEnVMj0YgiJOhoWN0OgdJ
EC48QUnD1rjGZEOF8c9ICnUyaINiXhNcQfhLXHxupquZ17M6MErGtP/zJ26211/P
mba/4iV/oufLQlXMwo3Vm8YctYh4r9g6jDAEoh04p28c/Hp3D5dyKwyvAsw21ONt
/Yg0w+O9Q7fXKOWSAqqlQrfG1WnSfe/wFdiQcqs/FeFHSPmULQ6+SVTNFS+XsCKD
ANb0mTRGVg7WcGGCsuDIvDhIh+jp4SFUWYBwjJ/ryoPF35Kv3AHXMYlfsJLy/krB
Kd/gEwS91bd+PGSWTrTeMqTRQs6P+qS57XIkZ7SzV9NE3e/jO7iYUUDnq8AQf1Jq
yBJ6p9tB8tMqb5qGusX6Gw8nNj3+HEb6Ls03T7OUjQW5utQzYPz3jgjZDyfMSUJ4
3fISmpDAQMDIeyTy4UBiAIo9JxcRmEaHwfdWmTDqiYPCa1/4Wi97EhVDBn4cC0Tt
m7r7+Jhiuo7tas/pdoqdQfjzp14QoJqIde1gowTpV1tMap2n1A8Bcx2TwIncu63y
Jk8Owgd9qsM1DbaySp89E0cuWW344zsTc3ObAmp5CUEt2LVi1I+YsWErEauwfLTu
Cvid0DEdV814SpEovUsBq8PvGnuBr4N5A3G5dulEW+4DljHiEulXHtyaObbRHWga
JETDYGWPRDVZ/83E0qHap+84oHjp5SzejDAdAjtGN8PnSiut+wVjKMeURgE4rD4/
hV5jlGoQ+bu5PoAlqMz6ykIGNXbRqcSBOuS4yNh6l3S5w+FUNzHOYZcWYqwnbqyD
vZUOWNw1zsScBQUMWMP0xwTz4u3UT6+4gi0h8KIvACMLFx2MPgqpjDZ6S1b84fI3
njNQmwZN68MoJii5iNFveI9BF6KidReDJC/1zmlThKuzyHbuF3/Vnnpwfw/6QQ9b
fTWyBfuVd0hCYDuaxyV30/kyJj8RAkoSNIT2AhBM1gRtmZVQ+P8Uk8I9F9fsXEPN
DfGqrIgLc5xeRc2iQbXiM6UGDalr1oo2qkllqHowQ/EXSKZp0KkcnBJQ8pOsIalq
oPvoMot2e+QouFzGsFaDc5i0QTsJWrOeQasfV2ytwhlGy2BKEaD6JxbDcbEP83/o
CZOf0YAH+6CSndQaL9rC2WvFj40vbaRD2m2xQ8HjH4K7CuJB3ap4e8HPB4e0pSd+
WwYZKX7W35YQBCc1XIWKWz2dJYhOqFjBowbLMAVVjtlcxteNL1k5S7WX9c4mf+RC
GtZJKzgu8BYyLaYFSJu991CCgUCezpvliqj5mAcFbYrnwZcx0Pzxuowi5mefPxAH
flg3GLKcAS4w7Q6OC28Fay5qz8y/Vn9VnZa1Jlgscm0P68Szf6kZzH3juVdByOoY
uhIfc2Ygs0hzwD/UDElzRyIs+q3b3Ne2pC8pwuSnNmRrmcLmadDGP+5BVud7oTFl
04zgQoB+LDG7a4a7HLC1HTpVXmdFOKaEVROsUc4Eed+h5hyYv80QpfIDUyDkhVDZ
teCMGf5c5JjpErPNEOu0OG53JCWgAKxcQz42wJ3GBRZxgicZx9SlxYJQw2s7UzYu
Egl5XO+y0ttL8AVB7SiGXAzHkWm4WTmICBQ/n6IkxmAyaNTQGr8kmj3kJSpflGTq
FKCzu3dzx9m85W4I9dOM5owQlN+TsHZQqtk35jpRf1cI8CFqSNKr/OWeS23aXcmF
ubRYMfEP1ZIzFwPtA6QuvuTc6N/32afpx2bhoRi85fMnw24PUFoiZgiTHVUJbjRN
TPKHKM6O+PVCzlpPJ1JeKf8l6pEEv/tSUIrrLI6svauoBOnDTemLbebtP5MjBpeb
VKOcBjoNOOYJC9ZQDFR96N09zXZmsWK+jUnjJZ5XSk2yKpTNPw3du+rVCQ0k1z+o
Fyta2RBsYaN33zwq/cj/ruc2ZWhHLwcSVjsA08+ztt4F+BiFqLWX/wxUgyihUaYv
fv6UpK4RJMCLJu+LM94P80+JM/Lw6EGaH4ey1/ZscdRP/TBPgS6Ncq22eyu/amX9
1XBISYSxJnlmuydm1qAg5/HYBFYwxi0Iqp/BUW9EKcEVuGgKFXWMm46snP+OF9q5
YaF4RFHLFEufqlw47Vwkl+yEZGvhHAvkxfKOsr0Ck1LhRh7p4mB1JaplFLGJhHmu
pjOHmzTUzk16PMBvOvd3MhWBlreYqBaQvO/SRjOZVh8pIwO0jGE15oY/mcWUG2K2
FG0XvSaISNfNBvaJgRIJ+EbLShjzDFJ68pg3vWRu5kEir5HeUkaOEvsIDODgRcuK
FaVT0guZ7SqfPsPNy/R8BDBFOWH59hjqfFQttrM6q4lgZ9G5xSy+kHe2n3hFEX0c
bbpQtWQDmVSabq7eeezky8q45RaXWos8kIqrsuyi9cUhXNB6FG5uCsZ3NRgFKcdK
XUt6FA3HqmBRr0N41JCu8hjerwlllZ44Cb0gm0PUE8pzsnm2rrdP6zdYSlZptf20
qjF8Cnkv18RWPelDthAIoVfU8WwTZ2RfA5c1ualTh8jmbdUI5l1dB75+Nu0UroT5
VI8owF3jmq87fuN1nted29HUNfSPsx5veMMRmdU3rzPdHFRARS6uRg2RGGRn5vL1
ibKubjHuIkUhWeJZxkIohaVhUsItja17E0nOwyaJqvpffsY6n6V1wl+jKREzYCHi
qQPBm3E/LMu2Pw+t7tlY/5SeRH40p3JkskT7w+q2yKifgVy0WWMqWOXaoc3UHr+s
a+qrZN0+JU+K+8HjnVRKMsRD7FlY/tAfbDaIZAfPsq50S8HrmtcfKwSRtduSC3Pd
dILhX4ohOyJLh94mkd6f2YfYbUXuwITe1R0wtLlK018X37hKeID9eFwvDei2Uozm
ahoKvCkxXDePbnStVS5v3KhW8KmZxQEm3uXgrBsCLrMjNf96N0Gaf56Fc2fxolTh
dhtq0HKdaxEObf//47FEDFXMQYlRUn2XaSXEYtsjp/ZcpKTAf/14K73nkPM4Q9sM
G2xGuvQJm1p6V0dgrTOYkDDNFTv3k9lXEyliQoawqq2jctzXYxuGHgBT3tMeDb5i
a/hicQVfikNH17O5bfDplEtMP1gVSiM84HSFMgNYI3Sxa+OjEex9x96zeghd8d4o
FvmZmsaFID1Q9tdqfmV+mJi7tg5AZlXPaCFFEhf2Qi/PXvplxJHnM8Yw7HmcXXi3
FoOwLNh8L6VnaopE+Ux6tmPGPU5EXxd/o+ddnwuNVDDPzK/pY92nwj69IM/nRyn2
ekSK9v87urPVKaZ48u/xbvnNO83+BxxKpDjmNi1H0ygWGKAxhIMlOTg6PfLN5nSg
XnN7GseKeG2htOPaqHR+x8X7x7iemm+AyyYaSulgim11HCElHNGxbyRhQrLJwstl
osLENRstNUEbjt0/Mj/o3snrXdwuHvM5SUXtDjjADmhmizCtFsEzxHUoLj6rM7yL
1diEeFOWQWigqPju6krVbaIDAhtTR4hc7E5VMpeL2hFGt9oZUtJP1tm6qfdIksvx
yjEmw+ULWDFte9JyIAsH1UM5nNZJ8UZYYcdcO9eyHDJ6H70g3GTWQtjf9hfanv9v
4ouE7uymTBinBkmQEcrOmt7DFPmKeUoc4gZkVR1CZ2Bl1iVQBQ2NnGEGLnlIXHVM
iT5WVA7FzV1gKkHfkErmhu4/ikiMMlh89RVgQuu00obCeKjDt4NJFrYisPcKPW4N
i3GAA02dwpYSHtx0jlcuXONaNX6nYTL50EuQHAWEKzG9xiKqzseAyGV61Dw1n1hK
YxHawGBb+Wb6D+2NlOaOEVzW5J413parNxLhDsQClgoOLp/3doxXqivzE14wtoy6
VGwIeEMldUJ3XKp/KGbJtU4VgojjKFfQhcYqH9G8t9J+xr3xt1HO8jZs8uvoehae
jQBFF510ZvpRCIGCIXeEaR0+/L3286Yr5cnA+AbvMhIuEYxqbI6XEd34V+ilfRKR
iR1kKfANd3IooVnK80eiSTF2EpBglvxJ0crhhQeJkqeb2CiA673ypcq3rNq1RyrV
ZfaCyqFYbG1CPrxRFNZ9O4ConKr81drdiMKEeotEHjt/MgjCStwv2zPWLJELLBq/
zfRY3fHQKc6IgxJ1lbw7krsw/XyoLAk952vuXgA6KGalB+S23U7yWDahnZ3iu+Xp
5GlXGSSQ6zX8VnU3Ukd/25CTQ4+oUBP9FAy15VCta295Gw9VYdeMwyKDshcr3QIM
CkJciShuTTLZpRZboVwR0Gv/FYgkUWztuQ9W3HR+67RlH4YXp8SqysbSe0nt7Izy
sRjRgXxv0CElZ92+o0Uk25XNxfWIgB1HJZXycemdL04RvwlJ1V7S/CE1Ywx95oue
gPhyy8SwINpIRAA57cGJMlljLAwK/e+582umJzKSYjJnxHq/ASUk2wf6yEdVoHgk
NeIb+67G5cqMfdmbU37HPW9IOIeJOJByWKrSQ6doxZ3kjqNle+5tFwXlQuBvw+nS
6KNtf73FPrgvC7qBRsPmFDz/nu6LfwXAn7DEJYg0FNMNQjgrrXQ/qIaVTKbcZ8BM
QZvzWbKxFg3gytAJsnI/7zS4HJWPFQeN8ZmeTR+6C1H1FSCgSGpGC96prB520ELv
F08ikKsBA0z7z2QoHAFNtrxYebPIKrtyWYJdsaeG8kgCjbNx6WJMlB4OgzrqQlxZ
FMKoK6hwzxrkTqb/mrdaFkbboPYF30vNMYMxY+0/Z4cQw/f8iAj8G+g2nmK7Wqrb
G1ic6uMTtaZDsP14Q1HuA6DOTTqVnHbGR/uBNTCfTw99L+ftmrHW95FJb3P9kBbk
12xs3HxdTPumq0k25xuuHSLHRX4vaYkpQGNRdogtFoz5+n1on1hxuAYzKYJmKlf4
vliRZ4AZ5wouNbpbytmEThCCDOv6qOBEslytFiNt675zXEHmTqhSe3jRFNpb1LbB
2uCmRgIqG6sv41dLe1oDofS1bIWHkz3HWBbFoA44WCqRVurSqZl5owzezVpH3LOs
fdzKjX4py66b9YdNePJnuX8SWqyEzbVbrbhWZglmYldKkt9YewIvpDMcCx+he0Fa
5BQbA+s2rHk3AuRrL74mbAVJ/s/jijnDN5QHvxj/RrHykoTqL0iczcIhLXrsq4n/
SUcgXOSkGmC9KFD4/vKnaF71dLak9iJWNOMfX7yyfo4qIY2l8pEnDcCEjSaiQeIp
E9xnVpY9AeXkZGwthF/6t5ICKPmZL045ONs+QUMEjHJtjdFuA1L+voZY8qJpbXuk
nIufC3c1OMSfSZQyNpNuzIM3VQs8/zTPgkHeoM4/P1JB1xC3H7/6OnKW3EFhRbq5
owgggVB8GLw36OmatTFZMgk1M6qfHGYS5zxhpnPyyQdLXw1vGSdkJvaX+CA7lrxB
YnUx6Unr14bdFGFzlr+NG6mcW2I4TR7eOs5b1RQ3eOJQwlCwGul8eryJVpNQkHyO
1ylX6QzOLhdiuha8IJQrHGuNrowaIsWrfD/p8rTY8ZI7nC82kX2Lb3BDNS59uQ8u
Pe9rxNkfQctwN41plv3SfbHzZNtavpulg67QqIxyNLAsEBUiWGRRe5kevIyB5le3
Wo+mTbJ6zWHyd/jWdfoCAaNV/5Q8btHlqTzOWbIxBi3Y1FrOPpcPuU+PwwlFrn+1
PBL2frDXy4glVGefO8gmdlNEAquz9HjLZGgj7aujyZSXFe1L9WShTgky2CBJyhSq
w+SVGAW8XLyxseCfwnZjeDgB62cjyD6Mb2KrtAqYs2xrtLZ7X1XfYhrVnPrmsidY
DZFUXeiy1tbUOyGei9NRoevzDt1xFtp/60EcC6rwtnbwdE/1QQqjYCOUUbG4vxcY
Vu6ktGLSVsiqtk7SA4TB2RKLOjwvTO2dC/qFUA8ZbGmn2GaNv4zDz7VsAMa+i0D0
t2pWG/X7wtJGE2+ymmQpSavcLXkzmJmBJOJ+xUOSriwdUIXQwMOFGG6Fwr91VYyQ
yehdV4mE1DZQ6uerC+/A/7S4jsJcAbgUgheToxadyRpZ+svGGsDxcjfraBuNYtuL
s1Ru1iNg4Vm+iX0xfgGcJLipqO2yDrWcfElWttZw2UxnCzlM7cQ1s6Eb+LshE092
lVKGeSJVeE/9onZgv85PoeAZhQCXW3CDUpfuciRBGjbcZCBvQLowzCCx/fPe1t3T
wI0FtZPPg23SrF1MOhMxbrWuCqcl8Pyi9JK+rV7TZxRmyAZhB8TEthYZ8tM7aofb
qvCmS1tQ8ZqCXu36h+VG5zYa4buWVkqkb2WnW2zlM0Fy4FYL+KMINhsy32jPl6Ck
mZMs+9P9QJGqiVgxfYxzEYqTOxIYvfSJqELYj6O7uS6/CtEO9fgQdBOueJOA33kS
prY1UWDym5Tpv/KMOFJGUUjQIuHNVIopLYS2568qpT8GKDUJEyaYaowaLeO68jp+
hK6/qsGqz8mRqBHpYjFRias9qK3LccJroqIULSqMRXV+RJM0onlQS3vjZpZ5xmWW
L84U+eBoy1wgRg3u/R5ff6PpzlhHycovPIz8xWRQ2MAgMCrsvCaIxEZCSdMkJZea
JPORNGzCnm6YC59jdm9cIxWRQyILDLg7b6PwVPzPr4LtwzHpHCnmVNcai3DHIkOq
d9e31rE3P0A46Afn2oKQ18xPmmXG0nN6rKl1oXa2AgVawJV6JK/qPmwy41mhfJ9t
Vsf1aiVql02GtIhNhOTIsfBv+VNzo2LKr6ivx084Vj/0xpwjKg6fgMKez34QviGG
/C9omn+cbNOV0sZOb0utqDGEiKPdwAXsBVecMzXbAyPVFaDeo5VNPWk58Caon1dq
76tYGqVUXV8VLuVtxE+PWKnIxOCaCmBa71zadzb4qv64VC72xk1Uk6uFSsBTrP3Q
C7LsQuyGhncHu7DPWWyMSJE7PRo3d51ZN5Hxo0sk+WIsjZlSbKADZI/AOPrPkvvg
bjaBwsKvKphSYi9YZBJ+bHBAeyKFuZc74OU1M/5OjyEcZjK8DWHZCK0+z89ikLbw
3ija4mQ/QWcqGA8Iy8X8BvwrJRqMo0v3LS3waZfOsTZX5mWGY422uLIddV5/VLWC
CaA4RusRShLuEkvX8kwYrpzhNhojIi9sQkm84EA/+qoDXFInojgm5pgNMiLjF8a4
s+8LhfBo2WujM9fHjE6z7N/XexrpjnBqiOEzmmE8LPHgM4ooFHLzlepniFNeDizR
Osh5Z9rvLDKrkUgK1Wy5OU92umAvHBTogxjvUwzVKlykLCBV69BE3AKUUC5zq7UY
Hu+8rc5Q6oOGvOtqPG951r04REgoaScSLQpdn7p8aQOFu0zFZYw/9JLU342UHaCT
2n7YXI3Hl+WpJUOrq6PAEGn4/fQWWOqY2I4cYSIAqkm18guP2BrD8MPxNa1Zxbxy
LFTL36BoqHeM+EygfgYCYP0B7ff8zkhQhBuzbF8mX+JxzTAGN06+JM08NJuOvc1y
7XZf8/QtxcbiXeK8RocJjr0x5JFiRqHrIotX9nvFenP244j2LMNupCdg7MsmXTqN
DYXBlJooNsVafMBzSCHIQIzBPhrc8tukODs1hGzQ690zkjAu3eH69mY3GU9ic0EL
nRCPKW05dIDh069FHczMY+O07d3FlIWXJJQG4gp+/96mdm+8b3cJgXaXHANVZTHk
vl7R+wa4O4pF3gmybX7zfXsu+qQzKmV4Gj0ZQ97TXimL7IbH9Jx5vVNwwtmoOxTc
XvZm3jC91Ows4oJY5CUgV70JfaArk7J9hlTBKSg1MeDhlIfevfN+FLDAK9Uwf9RR
bWz25UaWZMyBkg48doPkPRDvPq5Ke/0feffKOmvu0oZY07I1k1wp5ktiHpNth3jJ
bOsqKwPX8B231JNKWPggZXsdboiQhJAmvqbMBz/QBH95ajNG2N2O2agT44Y7fgOw
5ADFBJT/lTctZdulMo/T0B29MOOi2AGjFCqHcgPA2Ke6UYt05avTFnVjRms7tqYN
D/tqEe+JFDS/qVZxBd1UOHztGK6tC+UTCusx/bVm8gJCtvZLNPpDuU5Hft6lHvDK
9OufU4n8426xLiWhCy3r5PdSMDzPMP7NRqWWj4hzqDsFkdxfc2LD2HyfR+UxPiZp
jy8Zxn4g/NntkoYkA5zCoDq14KKdoKpaG1aPvKAldBvhwK3HHK/OOs17BBoi30AD
ZKcYQyzLcO7DLN3Dc9NvP+xpa0VZ/azPwiw+Vi+O8gYZ6whfMkTfXa+JJCcfs4Ee
bh3Wu8ezYPKmjzl4SxKI2071YiFhYi0EhDU2tvO+afr5vETpaqtRMziwaATKnOIA
IS9eu0gIcqzHR3UGF3d1urM/KnF6382gCb+myWddaqLX5YY0B1jqsr50Wj46umkm
tkfucgOC2gXuw3YUjLHaEyWmK8rm4eKVpjFI1iS/ga1GGQiGBH6v1p6jFzYrtx7W
Br4CUnrtBldS04qiw9RoOCikQaUoKP2hzxRiSnPmf0jyW23/tf6xzIOviPpdOWQW
S/of1Z6iHoGYBG5yz7vN6TreXe5mdX6lpvFF86Bl90++hlaUSJggiR9bCe8cvyQ9
V2J8eNPr7v+QDbjg/vUq6oYbjLevL0P4GhkrB6RvVukmr82sPGx/rQkiwAaFrFeg
9zXlHSdZp6UPxgqeLCAddv1WoEU1rhe6cnYWDl417s84qSjvy0CukrozI+dHFYgG
VJJBVHMqbjv13N5P81ZxjCVSXZVEANf9/8lLB1XMjtJcZK1VEFgTvCvnl8+KhhEZ
tTjx4E3aPRhvpJSG2J+HldZO82xnOYrJ6Q+9ow5zt1X3wZ4oq/aPbMtTlW4Xl/Zh
etVErQq9r10nHuMrIUnxi26USnnQ8Xi7+kH8euU2z2Zyh4NVAHXO3ZWuvrTYegL9
uTI5w0y8ckmi2nx/PYkuzFj0cOZ1TIMMaNT86oc+ZIZmIHgEWNW7VP8TiG12Qofu
+Vt/eZ64NXgdZRMB/K0tb8YoWiYsygSHAaPm86gAU59Cbf/YjYNRDDmXyrxBjtL+
ODNIW0jtz++NdmERx68p8R6ibwqW7V8jsC0aQxF045ynRJEJzvaAIHJ8p+o/t038
rFwtTx7XuKEfFW+0EKDAgHozcSAokkirCbpJzBZ8BJafs/ggHKgfVd1q26jyt11d
sfeplurNbdSIYEbkasUMb+LbzZRH+x6dN1R7sSIeV6DAN/WQhgCmdnBSJyrq+vUU
7Ih16dZ9/KFqj64zZ5piOBXFQczQUioydupx1Tqi5zNuOqARsmN5DqGbTixG2lNO
GIsI9fKGCB9HwaqwV90ccVpnquf1ru/l5EDXgvPf5iA9w45RWJqc63ibP68Zr9hw
OM+DDdYJ8LiUjRrq1aeWxyUSzHB4yV4cqWL4LHyIrLj5DydkGD4ILVirWyv4/c5Z
eZkQTA5srk77g0Zd9grdmfD3oPDkVwVHIpsdFs7aOczMsN4yowm+MjYWUT+h0PPh
2FPScXSQzMHgBjUxXJ7Se91I70w5uNeE/8jJx+YHiCj4lzDW/tuWhsP7JeLzC2ww
pq5+OOuT8gNLaPLgsB8Cl7/9Kms/2zDKyT0ugGhhDJ2r3H1W8RiS6cBXYZx5iUTX
T0dvhge9ICIh6UxQs1Re1Rb0DWQ/g6pQa5bQdIyJ8RvFTkrEKiR4LqLEb6Z/PVqb
tPytpqmrlShkP5RVr0pu5Zvb5fJoEDexK7/Mu5XWT6gxGCc3DV9J29xxtV/V7ihd
nyJQm3obfp+TTkQiHDzlhOUYs4IWT5uQ3HL8l8qSFPDKPwFn7PHWlK3r8hcGfV7H
D5v68BWTkdf+TyBvEwBzuZw/yuewR1NAklyRdiEecJTENSBJ8jpQCE3u/FHqCMaM
+NUX2W1MPTQcQZtzs1wtrluhY5mjb8MMg2lq2Nm7Q9hO7Xg0lEi2EjJmNTxKpirG
BmozpCGCI77lI3eEHtGYL5X5YItON62rY9qY2ewxCzXFyL/yJsNDU8TcUSrJsjmM
FIZ/BU9TCR/xXVA+6FTqKo/M6dckClFOOwg04OWXCVQ1sVcqYz790ecAwMr+B9j7
AdT2zCdWKmfpJcFjcdLptMO0dttLp9Zazd2gSONf0MjotfE//fyAJKnghibkBcwh
mcVa061E2SF82TdEwOX1FULjSjJ7fEYWvrTSxM8wpQXpyZhqWjBFVKbMnW2zdMoK
3t5wuy7G2KlzTyrhhhu+yrRhrRrOq/pVZ09ZChc2eFHhTyFp0pnSXNdmaTwzcX5Y
iO9CP5BGRAObCERtzvZcd4upGGwZS+LLl4lf1/i3gOOmi/0p/Byd8CP/GRDCnaBJ
C5XydXe4fJyI78/tpfqHrA286Xm5+UvzUsKtJtPF61ldNhZiwCqVEl3ft8CWAwxh
3YEu99c8Vc2DMoZXzTgJw8n/BeGTpCb93cmqRx3eb1CnaLKA95AtFsI+ZnI/R0vq
3rb/2BSiW9YqHcFArv4vzWiG4YzNChSvU2Cg1kxisxOZRBIl1o1055+Zrt/jYBtV
vjN8lmkfpTQejW6YtNtvWvln7EDg9avfrjYvHyCqq3XrC3GsEOLGx6LSMp3Q2Kpe
5sIP3K0E8UiFAD3PP8Tq5S2TTfmsp3/Yo0WhlM324uUsaZDlY096ezz0F+aVmBDC
kKtRsaekcyqzjEcA7bTcSTwOWc9ihAVAEslbQgCLUgX23la5KNPQ1UxSZkCVRyR9
HxRTjD5uVjPQRFG8g3cxGDf2jkg9jQqtyA732XXbFXFiLpjatwBumUUrdVI2JfIU
eG/kyW0PpWmVsfwZWvRxjUMXzvB2l1IMZgiAGFCyR6jpbZ+zsf7C24N5yXJh7oLm
6hSQTga/zaLapfq8iHEeYwl+2HVZ0nQcNVjjVcyUOa2CxB1LQHWozAh3ZmEpwA3Q
AuKFMFIGp/XEKu8H917v7GEyABEGmax/Scc4Rq/90WWVT0S9lrfYwPhpsJgcWD5L
bkMYNgYku25VxBYb1JKcqwOZzWMjHbxsV1BLn9xB9OXJBLAwju7iezG1B4q8EQwP
dUIDBVQBscWDNYQpTfT/PGLS9DAXtiYqBi3ogwqIr0P7JliZuUy0Dkh9CRPd7+C3
b9nL49vrTXK6VQAljQovA0AYFnW0QtGqxA6c/Opqk6PPfnyVAD8oMl8eMBhoJX5s
QXnOxGy8MoVvFeJCmT3NJ86CV0cYYHTFUUiebskPnORNg95K6U+qaPZWenVirMmb
phttDF4FXMcEbpMWiy2AHnfTds/LAHybx0Wi2YypfsjO6xDHSljqdk5lTiWlG4FD
u7ooimbAk7M5fOXcqHtrndjTRZUKsNejFoUNdq7k2Z+G9NpUtAnmClWAow6PLcML
SDH2uXtZnb6jaMrR2+pnkGiaCamD4smuuLDG5JkOh9m9+GeUDjv/D7bDfWcCCa9t
4ir/c8lnc3uvHZ/5tg2HLWXyf9mBn6BoqhbYf46EsEn6GNvMn2PyZkk03hvvV1WG
FwJTKH+NHIObRqWj/SHwfjbac+egKklZ6Brs1Q2VPvtF0vKBr8s4Y3+l1Y/lf4NM
JkN957AvfZyclfq0IwSeUcpBpJEzN8JM2vSXKfKSuC0Go1jiBg+PPmu5cUNrQF+4
kF9/HO8oYpto5LuTvVMKzOv7SUFITbBj8pII2CfHlgfxDpseBcYkaKl+SscEHmWg
HBvaYQUIxfT9mZyIdG8c58Ke3oD942+tbDddVcDkLYPlgSM/YD2KTnm2TVbz2yPI
yiQE65cLJ03/LgBgFj4tmV1V1JZkR+QJnFqUta05xX4oaHyFLQrhLhm1XgPY5cFN
8Dj/owpHSeNwc5U/Y2PtDL73Jkmu8dy+cToiMdr+4KsOTiLAtrL47L0sJAuuKXHE
dY7d385p2yPDQ21d/fMnLIkJUk3ZDpYUD13Yht4vKIFm5ZIXZQq20e4kbtRgqOEU
EeMExGIGn5T12c5qmwyL0kbKuel9dNZdcOjikExthjC5a+/yCbAoaEPfxehM2lgN
7Uw5Vu5B4/mQxwRdJ6w9TDejXf1RM+X9V2bO6g8NZvBUCmvcrT+2idvJNaV2yyVM
9w23ducJLuC8aZRS2fuAnlRNGLaPEzEKJchQHbycv1JWy2/LnF9REbwscKOoRutb
v7GrcnJIUxa93unnbWm7tg4djV7+GYQUz73jAzGn9oqZ1pRp+k+aBQpxq1Jdo3oo
Fkxzrb+KgtbZVZZHsXOw6CitF6L98tiWeYCY3tEoq0fkus3ZHk/oTH8iGdtuTE/k
60nJW37JIM60emd6I7otpaJfOsu/68+CD2VzrlWeujGh/pP1IHdYuHOKERrDENl4
fGvJV/QuZBExqO8VnHeHW7KkOugJWc3D+usv9KWIDr9k/piFvM3m4MetFbn8UPWy
KZmDKHCzfQydX/nnPiKQPAvJq6DXDsjj75ULXIpdl0NaE/9557l0ktqcIuWzvRo8
sIFIMzz+i8hZ0p7t7Rgj8pWMb+0mLJo9H1HBdCujplJBoepH+hdjHuNoDreNYpgR
wfk6KXZaWl6bmHgemZkx1+2+ldQ6KDSNaJMv2Mm9RXfmcRzZNds4SXcnBT9O9JGd
6hx5KPz7CNYmFpjahzQk3rX96321I6j2l7S+b59WN4Zcgj2qHvtbkXdnIIhW+Qtb
56EtSZFIl6lKB97l4w/0W7Oo8LCMeeUVDNORKi3aGPx3D5m7WjI91GRlkWVLhlU7
ybiCOWz4BHhbmHTviYpH+VvVztYx58oHsAImHg8zq3zGTzZtcakH+ej6gKyjMZkg
FU/ZXK7GNWicU7DXJpfMuNTS4BhVPbC0JYR3uL+fC4rLxvZTj5sl6tCIhfpgjRKo
jA2Fshg1WmTBw5DHT0qs8sEeR/qe7uP7Ml5zR3yIIY+nBEUEU3i3w/PuFsP7PaKU
/+D/uDm065OylIYKv56BbgWnjHaqIB+xQXvF5A2eDkZ1MXikkwt2ULw1Vcv+QKTT
mYO+uXQwlkNLglcnyCBMlMyEBAZuTcHuveCtvjCdFeg7p5ATxMSqsAuySbWSrU5q
OCv7Vqla1Lgmq9JJOdrknJVIjKlFeAXkzxI4JWwHm5kllEG06Rxq3vkJeUVOz+NM
HAg1U+bKli2fUsYWra2bYrhJbPk/QOEgmT8a+juNnEn+tUiI6paDyjVDfYWJZic9
K9jFrXwjz/gfpCBSctcnK2JTUF2Pnz1xrvDzDJNMpID7uDV5L9qHcjpkKRb7iWW4
0fguQbtoKdMFOiDXJLBAditnnEh8Qwe3z/hnYVXFQVaD0ia5Tgzi9gkgXriISl7I
l/pOt4ChjkZyVmd/dbJ9F48FNCaaBAfsRYp5VYkTP5rLUr2oanwcx/Famg+9jcgL
URoVeOMItv1RhxC6dSa8zD+cUTjGGbJUt3JAfo2RgLsl4QzEOKbM5JP6eXWFwlcF
MTV3ni1qsZSRXehNbHXSNfAyhve4jLw43y7ycQAdyUu47/MhzVwvMBBDvAtev4/x
xPUmQawl5EFq/2ByiSBed7Eb4qsPNzRn2PxeZ5f8oOcFpvOhpOm2gVAYONwiz9ul
a8SMzP3gOPrcFi5HObrsyuEzq0MDWH4dPrP+5+/TTDZIOC6VL4YZF5piIC8LzCqI
3fU5E926gQ5Dn7LxjZ5A+cgN3MRlZh/u8H26/zFLmJygm1cjZRZ1hdsyEVr9jtES
9bAZpZmXfqXMUEWyxD20d4duRt4lInnw7PtKd+phWWe2g4ImRygd1UxCBxs2FBS6
/o+cHrD+6PKw9O1joAqZSLIT1a1mxNq1HEmIn2WZ5WYLCYmC0QJskxDmUhUDAOGo
q8i5gFTD4RSMoHQNlonkU+/RchmwmvNjFh1KVeh+tmXJUj49vjnD+BNOCg4ebROK
mqpq/HN8u2f60sZDhMGTxaDKRKbTgKYxo+UmD+bSosn1VbVYQgzFaTPdGWXtNIf4
stEk7epiAmelkO7CRORk1+BVVZZPCOaJQi5HSWwXlPEBL6qWX/K6UL7f9E9v9VAQ
l9SP5XXrDgsqw077kVBFQXwtgJ9qUZqHmIH/ir2fXIJtx1rScCroY8FChk6hsRLQ
LFLRqKtaBR78qcNI1hMvmD6EnThriDMyCS3f9B794AzmxykQifS/PB/fnJTzVrrw
6Sw/xK42WVvSccOVEyi5wzZO4X6pqd8TkiTZcXgA3qQhFpK2bnAT2a/jTSFdWnmO
3+MADwXwm9f0bQGYZEFhPhyzCveuDkNjadEGsXSYTBXP4WS68qJuujHswmNEL/XD
KIePULnYDj/vHEroA6mRI6Qe/jFmPRO9WzvDHn8y5Mhdyz8bCw5BjKVjEeIa3aoo
dr4aY+grFPBeJfaEEo4h+Vm56vrofYUOOvIOBw7fC5cWJcmFErxbCXkeap/wg/FB
JE/fdsNmjI6K/6GPUnAiIN5v6p8Jsr9yZ6EgeV/K3cyXg/mmLi24HTEMQ6iEYQ03
5CUJcEdJCdzqaW6vyY6UfOKB+hWZZA68fOaam/PE+MOPYXRy3Gm9YzFblcnLWeSU
48A2sdZi8eB692zn7XyRB72IYYp1DhnBSWdC4/2g/vSrFaQUMQ8AAhRMzCS8n/JP
VzaX1zvCRSLYngFPIgybhbu0V5CHEOHX1gDhPdi9rQ7JLA6DBlxVpkwPvhN/5xZ6
A1ja3XjqCsoMcVOoq221R/cy44LUxhqYDKOLMvVrrl7W8cXSHm7GucYKygZz1a5Q
z2SGnYKlYnEMrGe8IM1ddu5GKtm8OBqNkqw/3979FuCr6j/qf9VZLEVogYbtIKHt
HjA8DUQXAsOOs3j8x3iauhgZfyT5OI60zPS8k+TMTPjNkSpsLgl4uJUvbdLao18I
laVknnK6IW+AQiAyvL17ZRIv7GY04YJLOMOUAT09mkzMM0of5DQF9YjMrmxEQUmP
BNTj8GAmVpPK3VpI2P8VTjzkCtN2nlLWNGIeEYKpauSUvPgwlKrBzIkLchUeFW5a
zwft6ZTWBv2TTc3tmqFQzID7iWGeTg6E1pAlwDWoIG5Iapg0llW8ORNaDKtAU8oQ
4E52NrCswlzbrzis/3o1hp6fsO3Wnwl/rQeadGUiS0tjbv3aUwJouTPmNUiIStWd
qMVcN5rPrNMlUYw79sT2X4Qb/IvTZ3oiZFg53KQLEob6BG2XK8pRsthvYP7TqUf7
8L/1EmH1PwJdqqyajI7FOWSO93EDLTWxs+U3DuzboL5ULXdD60D/mB3Usu0/ciqF
Z2kUXo0mcj6DGWm0XEhR7uEwItLU3L9XXMyTB3k/wUmF7PFA3ukHeej8pVsGcmxK
tLPxp1KN1ZJhhk4cUbjwZhs0h7vlOq5tIfaEmWvyjY6LwI4F/cOGbaDpJmGyApu8
Wo7WTO/PHm+yKI2XXXecTLXFdIWZAahapdnqw5UOF0VPAe28pXDB81okWBTgd5qA
xZjMC7ETkYlxL2kVPSvKFWv5pTVZgUjdU7lvHW7Ephh7JMZDaaOCRv7Dht1U3G5l
2xUQP1/ORi+57GcJZTemcwxdni8UAYLrwdm89QxWItiQQDmbLxd34topgwlLuG9f
xI8HsQKa12GWfozwpdPX2bYuPX1U+00lfxJTO+t88djC/7J8D5Ain0T8bomZWJLq
HLHKMW9GMasaFyVGMpwC0T9V43wfKfxl/fBqQjeGGlo8lIhC8lbbdI2BmxWQ3nEe
+RIgaokaLlPPfKynAN7cLGxb/adIasYrc3M4xWztfZUmeAruXplVVSjOnaie1p55
oJwX0v8yqctm8ZWuiIeD7mwyM+SKb36f2L9uQg/dIwpPtfqQQq94Pdu8Xf+zCmOv
x1xaknZ+XLp67zpkMbOFCUFnmbYHGzgXnkJEMMvjwfmNw2pbZMDSg+PbuD8HIdLg
PFnTTl8YICNnzGtv87P750cE7apPy8n/m5O9GZexqOziXCPnwkdD+6h1TOPhmrS3
1MS9U+DZw+YOYxJiGwMnvhO+OOjahH3i6KF2Ekh7rG/3PoDTTy7z8mqqa2X/sIkr
OHAeODB92nY00d62r4LiX5bHQkwgjBvdBAr1sxwryLZT7KwbV8RZeiVs99s0s2m9
vPKFTrQi9+qCHs9QVQ8bIVrzj/4q+uLRsS9GXzo9UBPUacRUFfp+WdZ4XzYwd2g/
lEBrK+wpB9mHmNmkosG2t8EbdpUMwSsHsvoSSXmr3O0Lisl4KItCjNwpehhw2B8F
sjWOEX8LR4dEP9Jmdk9EyiWJpdFtsWrNzbM907QzHNrWra7OoQN9IeteJ6I3rej4
reeVCsccSCteH7ZXVPrJ2deZbkOXwEE4iTrjmXe/tOVRySShLyf4IbVqFouax8RR
kHBDMum4GPVJeTtA8coujXgyucVAgkZ2QKQshiMeMg76OL0VpCFXBSCOCrRNF6yM
bEQvcf/5s2mr3D9v6ZWunfJe5UBixwXCAq7IgOmSSxrmurEHcwM2lLDjFEWvnBLT
cD5ImGAXrz+GBgW4PVf+AokFlYwdRpTEE9bBslX/MHF/HHu2oT0D/PiK8nzYJ2SK
eOT/CYvoNaD2slKkeq/CZObDIMZxmohxjXceftvWCs1ataZMvDpftY4zbDxdsuwg
OzsdsYcKcB63qyL8MV5jmFFIS5zSpu0mQzv47pOciCkwSY23UW3VGCUDkU47ccvL
SCDsyJUa9vNB5Apu9DG/WA0Sx8EH4d9ynay21pi3bqi0uvvVJO35kMSf+DyUX5/I
KIz6W+975cUVSHQ6/Qc0+TuFi8RWP3s78ptKNyA6Odx+/0/kpFzJXLsUbCfbjyh0
AFXlEKyCttaIlIykoUU3rrx5sUiHvPhK8njuWM4Ht0zDRHdQjd6+BeuNwuPui3fr
ua1/8dx9oxpdXU0Nl/QQ4N33cUVz6+vcgLJIPU0Hq8GTVDFEi64XLXZXO3dlf2dv
YwkcapiJwPPE+/xR93F9oZoITmSuPvnSRhe9gJ3JYFYILAK8scOGAhfccSj31Vl7
ezlPGXxoo7Ir220w1XYd1dBTgtJGwvsJnMzxhEahNVPCGI0rEeqflVD2ZqWQw0ca
/cqMaFdHmqVlZrLe8aynAItBGtzcA/U3keb/C2ipk8wThu0e6QUD0Odo1e+6AL+1
93EUnzdEC/Zx61dghJ/iYrP2Vx//UQtsb049IeDEIFYiG5DhVACHGM9yfS/1lKTS
Z5Vs8LhyToAuT5QXNdMNEpiUAzyBZzingaMqKMFzZAQO3eV+S99rjMt1V0s5TA8A
NdjV7UdLTQYjsu41rj5xs2l5GcPHYo0jOJ0eeaQ/sCtZ/BiZisjyS3/vb5WtDJJL
EobifyQ0hj19fhejXsXqgab83vf/bXxOcNVKHzbPD2fDnUZFAe/LYhemeFJpRwDo
Rx1X/o7FUZTTKbsR/s2JD7tF0O/y1cpCcOXKZNux33zWVeEKYsHnmjqb+HATh/TL
YO/PQNEP69ovWmZM3AMDKwZawF5XzQBzQTYhADNLfkwYZ4iJWkNOUoTHIdkx6OV+
Oq3aYLO9EuaUN71uvy+V/EH9ta6O8ElpKNuWUGLxPrraeLu6yDa3Del/zfcHYBtE
2Fo3yKqGPP+u0xpDBe2lI+EPTmK/YM8vP6x717QYrUgEnJ7mGjEwY3D3exXK3JsU
0RFLiNYcqNZk1ce6+hniaao42qM035q6+ApFbWeT5DebG+1OO/UYLB+Bc+j+cjpB
k6UwbJJ4U4+NzpbZaCgZ7WRyrfe5xcYJ8PIQZlfLySpK8bCCtXt9IVKwUAxONeB/
EMkENiREk2qjhVAkVasydKAMXYN0syy4PjfCunc4FddiU5Etgk54sKUT8nAT9LU5
5XCyMiJDSPWM5k6GN2vFFGZ5Uw9RoOM9Lj3TSYVv5oCUfLZEQf91jLjgJ32DX0PJ
hvyDM0yXNqk9Kb2p3Q0dYObOWUsI823SZA2XkgkMCtK8KSUXeksjzoEmQ1E14EDE
WPOH+nEddIgqnVi3/+IKfIMKc3jlLB2eUYjr9n7saCHXRwvRJPUpG0uFgdkxGxbC
9im3hn7GqVtssxTDdLPUJKAfH/pql1rCfc2wZAJDpzyKy+xPHNZts8THpc+DIJOS
Kz5hj14zAXT+GhBa1UqvE1EmRltighMgw4V2PrJoXi/U1qw6bQBMAlXVDqQA1Q8N
CAdUwePwxyxidq1sgz/IjjckjcG59nKOI+YI7I7ZT2kpmyw5EFRNbCUCWt8YlEoi
7puuEVDp7AhTfM1q669FWzs7aR9DFoxzY6OiX5Zw05rk781Rzpbz7h9Hx3Ard9kc
M1uDCbjtHxLY6s7ZYSCJxZ0tFPTDiNehn/KsHlgZTMDRiaOgm+cyKZUdTXZ0itVq
hAeO+mW3/9SHxauJUUSPAgykXz4l1oJuOwUgSxg7g1kGOU92J8IW/wFEuBaupu4h
1P4B0ahMiVlBZoFOPtBSVBxNFB1vqbZPt2zViT2c7rKJB2+r84uEPTSgK1B3xMvd
DlzjP3QQsCG3+4LhZULD85JDhF0QAeEpV0C60lzPlE316+EFebcowIPPlYa8kABA
zzEAFZsG0FYL16XMvckX6SXd+7UPAoY44WE1d9i6EuM+mMVy5iGK/gw6blF9dg3n
TGgPzw5udc1rKHlgK/Wxq0dywZI+FVg/xRWRIr7xIBtxIrt9qYk1Hu+UtnIGLInq
GvJ8Dw8+i3/eQ2TeVDyY15QNxbweR0CLFghTA6aSu9ve9hvZ/kA8lx9dOpimyC66
xmPAh9GQ5UxMWbCfBdSl0gEQl/2sMpBLUzE4SrP0MRwiRAAUiQWzmrs1i6KLejkT
/q3kcGdG14E4cH7C4K3YSM9cyB4V6E9wjEmZMnPPDIQ/DNWBVQNmqfAx52DqM+43
sTgf5kSAheOB4U8dik7h9YM1DRc8u1R/8byNenlCoeyUrRh/mIMlpYB62jH504Nj
bBwpRt1viIKPNtxW7y2Srv/AOj7wEOiBau3vbJc8Rn7zpNbELMaBQawJEvVBQl4q
S1WAd1kRlMbfWRevmNnUB8vY/WSL3tHwPgNIds3edCKTVhjl731rPMsQ4O7K1Yc6
9jdFIyOPPQXuMJAyOkxqR7A2hfuIeDbotT+5Rca63+dQEfAdpv7LdbSg0rZAo/Rh
EhPjpg+6OWPvZ12JhS+izNH4wKybX/QJlBFvJylnu2quF6x2BQQLI+w4lAbtziZh
d8Fpx46wS2gT03ciKzy4hBKPNCuXammyktllKhIolqnaCe6FKsYE6jMWXovc9hpo
9m6RrVkc44z3FE7IpzChxWytXfsztFr+3oof/4kjrwdw6akXaGZ96FhlrOquyqCZ
10rBcfylIFRcvkfrXVSvIikaCusilEpDK4iOovaI70M9GkcF/E1sk5IPDgCpRcUi
OarE15z7EFV+8kvnqpiqP2i7kf6gNMzObOcA7bnCWEPKay+TxRa4pKQqyzWotbbM
+ag17kLGvcR/S3DqQ0b8A/iRFZcP+xmlXHVKKsI1Nl9orQxmh+8ZxZytts5ASgvb
qcDZrYvuWFeGxWI+ISKDBniju7FG9ARtAAZxzUIF2sJDKBfvHQ7z7evAL/rgvJyV
rFjKyHSj6QKqQmjDkR+J5X+z8WkG77InlrSQCcoTG+zN6vxp7DljwBiJKStCY/yf
RL3ORI5ZxCosPmRRPT5d3n7m9pk+vBd00z917otMqVEwVD/Q2UnClrKSIW42bhwO
GN8An4kX4Wtwv4QUVwN/DGMcAFqhvfRXuDBKpkgSzYcZ2CghMGQg3v1Ix1BOBFtw
fnSQBqqZwu1QO6mwXHXEsMkip9B3ud7VvzSd2VBWPHq3tkFPNabt+VnzPSSu1f2W
hXdHI/OXX8LsUMDWxC0iFvaxiWLboHBOgWkmPBkUIsfoNi2yFOgEiYU3kCX5QtsH
oV9oa0Uqp3ppxEL0zvCpjs/bWdGl8aa3G+5nT2khcUkMpxSa+TwVGBJHD+iDLrPb
/px0b62t6a4RJ3jiTtOX/js3rLzO2fpJSqpIR9y+t5uNMWkw2F9RCAwvLcyS/kX+
Jp3ulVOHF45KmfJULVuhQ0I4CjUUdPWpAgomdOd7BtCO7y+jwDSAAm7XchLcxlc6
nfkraRLwUZeLf8NnJ1XPmrchJl7Z+UL5vzlw5z376b+Du3l3Tm8tQi5VcaVMhkTo
cOhH7jpfn25iKH+bwyRu4XDHIyOKt5jGDtcKxuDE7+FZjLibjtIwQLC1uDQqcs2z
occww6a66M6YzkGm2u9m8lo/wWtmjKPyJP3vCJI+inY8TkNR4FvhcpkNpcaEVuUs
bqOWqt7TDjxeu0+lCQhlIVweYxPM2rdLpPWBEYiCuN2TUU6wGZT8kKPYEkAw0RKi
ECo9BAfoEREZiqhVO+zGYaAvBswt8yXddC8DSPvHcHIe4wB4poF4dfvwiwfXjR8c
g57BJgwiOG8QNTsemQ8xtrFb/4bVdDSukIjNdV3Vcg4qXPkKqcsRQwwfPUrVdndj
VvDWZbhvUIiZ2uxO8Qetn1Z+g0QUVMOK/Odv8lXb/FmMRzk6KAVFd76mR+vZ+RLF
ylq+tHwRtNaLC0KNarCeCTbTyqED2hpxmmDmhB8Wp9A5Rtriv11i+9a7GJ5269Ih
mObhD4mY25cHejqNK5maC2avZti+kkR8twpAG8NEKsChKiKXT0g2g+jpBW3k1sYg
3TqUI0frQMb+5jWIOUuIC34hraBAGVmVEN00GRWDWqkDYSNusD7LhqWKxzCGY+ch
YyFlQnY10mxoRIL08oTsqk6adEr+7sWenysL6JF/L0jAzZ/4gqSiF2TOdz5wXuaB
cT/uihmxzzc627anjMIUaiLIee4A6NIhvuH5OIUZ+NkNG7xkbW1HSIJoVL4k9kYV
QGuQS9eVOXZ+wmwGZQAt0ZctAVkuKRsqw6arsZgIKDwQvbQz26+o1mNfkRw6ksZ2
4DRGi3XzMCPtONsKs6IYPONQHNQgHoXrk6t/RujWZxjUO9U7s+smrbkeozw1xwLW
dPaPt9QHBnmI9HC2SpBYnt2liAX+xYtpoqyCkkBiFIc5o3QmfYhD3Fm3X7lKWvuy
LA/IHO5tN2/TtoZvyxqu1qEmyZKqnLCJEedM3wgzBZTwsVCbMZvM53BJTdQZ/G+i
/Hnuht5hbco+540Vel3Rmdi2xngdZ0dS8mydvLH5BaOyLn0g29DIZglECZbgYzrz
ZzhoaxeLy11uo3zBL5v6vLuZdFpG2JgwzcJfMMOPadnBqh+w8kJA+bgMfyAtSXbi
H4rKoS4DsNXkY+6qmyHkx4nCCt0kbQ+rL4Noshum2mWH1wNIA8xuRq3uzCGq/bAB
6HE8I+prwg2YxIZJAY/R2tGLM//nZ6OLD7JfYqYryqszdJzW/0ANQM39Bgd+4bR4
kD/Ukd9Bf2oNzKYheSae2AlwZs8zTEp71QEWPVtboNB72LDk7j112mtn2+xPcct2
/KI0EmHQCFJljNGzTn71atnuEQyQQ0zf2UaulCotWIGssA8zx/B41DA2kLliLT/3
jjz6MBd2cwdvLxPJVFk39qTxjDKjCI+ugN6fiIqnPjH/rJADuT0JtcCR3gpS0fhl
XJsHD3tE6VHhm7fUS0HOk5G2RiTkuqmszPl7ZCoXjvs2zbHKc3lbKKR3JwXUqpu0
Z9HZInZ+veRaQ3tTj4RtDy5BcamtHMEFmDRzEKE28m7X93pX/UDmzwxP0BGxA00p
qaGp8Af7K0aHY44rY3bEVRL1xWqPH3Bi1SANwY3WErpl4zZ/72KICeL5Y+ZYtBlH
5CbREFqcFtMKhopbRJFmx4xlbMNjDfK8T0g5abPa4ITDNIW8vFdXjgT2a4GTHTv0
nUwny/CpbqScFgR3DkBTezEMosFgcK8EDqH9igrLiLmZpYK89G8jCD//ClmHD3CR
zmkBimP7EaeKrOgOe+4mm+tx4i/rpeark9S/HvtBBC13CujK/Q2lhlN1Ts5ajJWm
tHIoe1j42rXtKdGWz59vceP9ynJEkx1TpQDZiqCrm/tKjGGLlMNBXhE0/nqueDSn
/mNSgKEq3xYzAR9YyfZ/hQ8yMq9vJB6fUOoyySeYcjZiAK+dLt8wtofl3PoMzEBE
y1HGcDFE6NEywYC7Uq3Zd+DEeN5XpIypRaKVLgyZTagPBf1fS6A0gxxkXMcMXb2A
pZT11LvMu/yESvl7tX4yjnCD+WGM1kKJLnSKX896bkdTK7tATxxyht6jztMDv+IQ
dyuQoRCXbSQtVyQ9jDiFwsVvvDyJh94GVIB5mjths5eKkLpyBMmtaXWIycAuA2Kz
zQ4wiVMAyy994K0rjzUeIpkXTAVSRZ1IJuwLuXHmE4TS4TT1NzwMPm+D92Tw3tFx
0+qyEgavrVTm3bqzXi3M2k+b+tzhx74mb+vlm8aXK0whi8FqFBSQR1Cmr9wV325t
XDOFuROMPe9IixebeQI8db7nBMKUFdf0FT6GfqlsJW4WVURgvZwMoSlgRMAx5Ccf
uZBVNbtYP1l+XDze85DY2SAzhk/0iv5yS9kecPMRLOmaPc9vYMTo+Sg2Zl/XKMko
/I/OevkN5Vg60eB/rZ2PlBKOrD2+zoKyJcS/Bj1gGx+tN+s+1TszeJFI8VoD1TLZ
AHNmQ1R8xzm7zBaIOJU1Rv/BOd9OCfUDDDWTMnl89rwJzQfwNmZsZuHOPJN7S5uG
RxAJ1HBYBIgWC/GRAHnwFBOqBWUaxNaM5ljFu2JQR0zpcZyU/BTAxxpx8JPIMCQC
Fb6Uplt1H3vExWc8/8+WorM7K/28kJvR8BZEDqIsIn6JQPZXdhBzDqOpBrYWoUwb
Bam8OJd6cTH++lMPQYiQq1nY6vv2/skwriU4/UOytXRQC1JwM8k3Fg7Wbe0N/3+A
CptMU14pqKXvRUnyBLUhlH0S/183nkpxCnhjhAw2QeQrDJmhNn9OD/w9Gx+jjDGp
+cRl5bzVAthmCNjkTMQ8qTUGxPBZSH81Mz3QJbYPm+eZBqHpLnArNSOhr1g1afF8
uOFEx17B2jePKDsA3VkaPxELf6Wr0yy5hhen3gtXUAYT1fxhe1yN6PovHx4pAlHo
ch7eK8iAcxXHgumvEq3UJjGms4KYPjJtodst6scWyx5ztPnmV1TOWmNcdnRIUHdg
tB37iXU0/S659Kg4R8qb450RXApNKQqqSNas/qsrSgzgTL7Z/CGSGwKbqXC5AUuL
u27nszSfiO2O+NXKIBW8uDFZuWqQtmY3RYMd/kwNCAZoV2VN/T0D2+nlaEVV140j
AjmzKU4VBns6f2HJDKOqV151D8ZNWqjkY2Gf2926qv5qvUmpaaPWgmGehXDXAGF+
mF3yrpgIec9lQ9AadfYfGaRsPxaXiBBNtzUyYLUtpXsymN5UegMNjvyWly5vyAbc
scg3+vgbY694Ky54r0d+GKtBLLwArNudjcVp58wVzb5sT7F5jEJaFoqKTAIcBkf7
rP/Fo8ZGcd/DWOzBbasS+kF3uNrO6FIahm4B4KqXBh0O/h+zu7UZ0mEfnxNiBcoA
owctnLcqOXwuYLU9ohtEc6JtpEncTfpuzeAq+YRy2SWAomjhRzWAImP5xynuON+D
+VOLn22AYiQbb+gBqOSJRGzk6/lH+MdTrLl95b/L8QKacBc+wybimbY8Flj90b5c
GOku2zXeCMA/s/Z/oE5oUo6uzupnXqUhd8w+dHcAke7NHwnvamUAS3/gz6Jjx7K2
6O4MRUzOdYCAT466kmqJKO4KalNWYA98uKIcT3KAG00z9K9AHFOTdJlaM+iEn4Yh
BbMMIe5lCtI9qiBk42ZNVTN6aV3Go41JExSjEFw3KXrzVoyec52/2n5+WQQ7Wx4z
K7A7fbdux9BxfmIUTOtCg5ossf3CzvuoTh136RzC17LJ8t55XQmul53GRW1VcuM0
YTo1TTzzw1ikk4Z5LQrSSsf+JZvvf7BzsTol2a+slI6XHR6cze/Yxw9Ydv2zAHC/
HONJg85QKpaVR1fjwR6WKDYWR5imQgGb8Qgai+Aq/wW6hjQJnpRSqn0UDfWA13NF
cRdt2TPO5jUE9tv08qmFMwE3ep+ofLlfTahjaE7Q2ZGQor7bi/SapFN9MtxeAKtl
ruHxYz4rdgxDt8UZv0NKGdCba1lPJk9SXmZwiwLeeZTR9NVgVn/9r7JjqAgjkArJ
HPztMAU5xCAVd//yyrNfBXL4RtwuJTtf3/OYdIvYZRjvSR+x6Dlu7qtY0F/lz8jj
zmfJ82DmVt9pQGGjMvRDreqwuArylRMqkweN8FQffrWyb5VBdvl5+Qf7DJ5RphYo
v4vMwxPdk1NUXeFtd0G3HN2G01vTFUzh63oRC78TQsGm2JK6gt9At/dwU2m39urk
hPZ2UCFert5ljGjF6FkNELE7G1akoOOYlPHqn1w8m5h3kyRN9g5Ti0cbQY/+PEQQ
U5oWh4KLPBjfLiNCexmhjZJI9nqYIqucGT7FQT9gqgSMIEr+Vd0X5Of8F/YCykXD
HxrNpPOaGZ1WLVxzSQaiPLQD0gSC6+h2sfU2aZc9Jjx6MHycDwMQxn/MxgA3Rt39
mP/hKYBijrQx/+KvQiEa1i9RJdp2f31AgtcobctqQT+eCee3W2U0+TDEVloz22nL
HRiM/hyofpt77lp+xbWUOiY7IHs6u8YFySaUVueioMz/pjFvD2ZdPQ5GcF/KUjfr
tLexzniV11Xsx1JuO7O2LX5lHJXDgALqK/eL2cnFmvwRV77/MatSvYViDvZ5HzzW
FAVw3XoeEpAXpIvNQUKJpreFeOeCLaVD1i/V66PJwiXyqIazQ/tneCBnvjlOTlOf
mDHJWYjqkXXjKBZ0O8sD8gnHz3YjXuY8xOJPmhXt1nu6ryYYxsr8y+kB/VFjxxTq
E0FK078cx9rvtO6Sy1R1ENHDZL8uThKzpksj17MXkb1D9yuPikG3CrQrnrsKhT1Y
Ragh5vIqenHwCs6scFqytB89e9VB2Kly6YMmEmczh5AidvzstZsPLtMGx4Bd56Ma
9GoaOaKKPndH7Y/ncGWa6y/3U+aARzR3dI2/2T1QI6Amh5SrF1kcVQrx60997ict
lgJrz/CEheT2r89H1fIJc9NRsMJY324wy6RuLTQ4Zrk5zc5P/hYz9KPRGhBCgYTf
WgQq5T1u9UWL9T+mverKjelbuJAk/4op+MfH6BL2RcPdcFTZe4FEPqBaTXjHPF6y
7Ut41PSz8Ta4zQz7oEKbLSs9Rak4SRieKp7crg6FC7bD4vckMi7LDXsoLGgW3D8a
OoxzO39m6HEnx7XP2M85SeeWHLE2rqfpAYldoitfxzs2sJYhbN+BGq63mHMYSdT+
lL9+DHPJthgZCJ0vJIg8O+QQxwscXbMqKoycGOu6/t/vjqPTKGbnrcJ8m90RkuF/
77rV6K5+CixtsSwEM/2XFBzma3QjUxNYqWts2s1npqFeC15S79WtyPS5ilmyJbg2
BiQ3+Xq+JPhZyrmD5dqE3gi9nbCbQHxrDgtwOV6qau0BhmgfgbZsduiRwmD9e2zh
lWt70oOX8FATGU19QMqZIoq3rhGIcF97TlUE0x9/Ms3J3ByCxNDbrG88nRzzUQIW
wINot2uC691Aad3u7HkHf6Zo/US6hkN+vpmtD8O5/s6i097yblYQohB6UqNQVxpH
/V/ZNdH+scxQkHmT2y+TgAHHBZH4TPs59qxQpAa/nMTnfn942PwlWDtOlq4nnk8d
jJss4V+jKnZZcp91RyqM4oKbPsQHmsV+t7DESMnGEuc5SZ5M724kLYlLqvtAWJmp
SwwUIA4+gJoZDpl0Olq5wgLI2kv8EuI1BaBQDq2UwWCYsoSHyV6RZWLI0bZ3C/lt
fgWDVc/C+xJQIRx9FzNRvNu3r+N0bKskkJc7OTXBv6MZ+/GBaRyuKWuuJ6dv06Ek
f6vojNZbX3pAKXyo0V/G+elsZGn7bEpJcgbpR6C69h/YAq3yjN0sFWYf1pXIyHe2
GlNg7eKj7JmfmDMFP1GeRIf5Hw/s/SjCrS43oxrw7E5l22oCdwnwI2h1YvsRpVw9
Qa8593JA71ygmUPqzFOJjOL/VM61+eynKq/A4VGqfJXv7ZJUjXOeR7M0VW7aUFHZ
pqVIq8Ggf37TJSgRcrIK3cyRP22zMpIVV3cXqP3YHc80P88j9cqT4YaZpLODjLxg
EC1P+v5/gcKA7yIAJhPdbn2u21afiPQk1MgsVyp5Al1ds67W9vWGUohS0DLG+t+K
amQ9W4D6zOkh6DeDqPO2iZEB/Z3i0zz+qZyD1xjOG+R7GQ///quK9yG/6HjCcvIi
YXFNL/73+4uSW3DQNZ4gBrPP2RYQdSY8iTaSsTG8fq0f03/NdoyLou+0JEdcwEX5
yycCMLuMLrLAg4LjNzFcZt17iAtlNK+flUCSKurAVuFYPdh7/s9hQ/Kd3p2hUXqp
ksAtDmwqrhNodkwoRsecxmwpFN1GosKqImI0rrrtpe/O7GY6IzuqnjlZ8RjlWxxY
++filWHi1B/9qCDzLkl/NB6nREnWrfQLXJjngfIZEzA4QUz/Q+86ToFGkc2lSNfD
Spq8Q5gqS4K65l21eaCJ3UdJ0vz/e7cnAWLfAfuSSOp4CbLmDufmf9UAOFx3dvA8
pgo/cDJpx0YdfL0G83DE8szsL1p+D8aFGMa2A891DNuPaRV2QhfsqxeaEzdcm+PB
yU1AnFLjg3NzsB/HNm2zjk6vjw5u9ieBloOn2Y1hIMx7mfDftSrAEmMD35z/K6/D
Y9H1zx6zSF6khWcD4bCdD40AEsZIrgCw4IGRiu9/TiLviPZkmVbrxH0eQsMdxtCM
0g1mG5qy9DZiFhA48l1DHRKNBtHlxW6Hhyci1/N/bmKm/LKFCAS0O9rKJl2Bw8l0
RrktATJX5oxQOfuYMHhwB/Wl95+HbVeRLjwoPsTXzEzMxb57mTGonbhDeFMye3s3
3JxdR/AoRMQ8bK5w7LODZn/faws67sZSYqlBlTxl/WFb3pg+EFZbEP89TBk/BMHv
1YToehYrkazuU0g9WkB7Lre8wqe1nBMStpIUe2X4o6OseSRuzcYYcjkQk8NBsRJk
Uw9gPSVOHbYsYr63IdrFyvFQpXRenbQSa3y8dbnlbvSkX1rETCP87xp3yqBjlp+l
GSATqlPntTsSQ/z57vS7aOb+DDsawV5LPmbRPfNRzU9XCfkywTUHQAj7tQbtBEe7
R6m0R+taOiCcwA/Bo2joIJm3nuaXVUrOYkNM2uu/5gfWiEbqnL1X84Z7iOp3kiko
av0sCQbwAwMERKEFt13VAG5m3WqFZoCsrVl3d22+A3zxh27aYnipOVfn6EEQi1nS
XzukzXu9KTJSfHWxhDtvw2I5x4pqCtvHvisg0sXbpWLd1WB/q2SM9ymAgj6l2Z5y
i7EcUfHcPYp8n/CW1H5lrjZK89EXTtBz6OZdh9JtbaaLOyxAYAhpNvEIOVqz568g
Pf3XEsJ8jQhW3/wyuXooGRqMWYBjT4TVtL2+vThDqqH3RNvUhnMJX5Qc0X6mXKyr
SSzvtGbfSjGPZP7TUvA8AbaAksqpCwCVy2+qqR0OKU8PZGGJI/1lFoxauGlu2E5l
prufPB8hGqyBQHf0BNfd9/8gUL4oA8n2N9KSW53U4Ep6o+PbUrtiiQfGgkgjEZ6w
APb2aLt+Q1zGaNe8I4HHW8YcAre6LPzFa2x/cLv/RV1Visi+fM5C0chBxlxgN3pT
+xiKUbZRfAGRR0Wup/OI2F/BpHbdE3mmfAvUqxAVTnlkuZiAutUikk4hme++I5l6
L+QZ5pa6/f+bhOAB88pQ/2H8cfe5gBev+uA+oEu/AGXuFjvx8rII69gwa5nMB5/h
IA82idGz0eqWT+Fw4eQ/M9Oa3NmEEVxDqIIXIWjI2FWJLKgK8/vr4gx93kNdFcnM
4u44MWJMt9DZhW0+5osvm3rTX3aMZU3bYXFPi8r7YeqmrkPBBA/DkuUSektpyc0l
yhk2SBvo9BbakTJxCT65SFbU45UWZGf7GqnBncH9gO6f7se45stSvR85tymi5XUm
mCX43LzblwY1LMABFyvhYJJw2HwJFMfGboyUAeUwWRvyQpn+0TMeH3x1hl0wmwdf
n7hhw4ONIITvD+AM+BkbTU5t2VF75BamFrJX9rGXaMTYSkB/G3sEaRA2HH+90HBs
DVe8IughE6P9tIoq3lDspkTL0etZoi2X8QlagqFuAzT7R2MBlfhqakkRxdOXcAXV
wFyJAVn/94bQhYs47ZSk8r3Ky7425rbH9owTpwEr3j1LsIGXmaaNwQ4xomUK0pI1
C5T/HRviVE8VatetZyK965WAMPihyep6RTA/NNi8LbEorPTx504kXnTdok3kIq3w
LSZOBt8yKtx22lT8WXjFvosFhYiA2AZAO/1U8b2RFZg981Viy8qBjOp8FUKHFAD7
/Unn/FU4yzKNOqwC/XOnLbbMjSyzwszpYcJszlPtxHAEOS9SeZRqTJql4bgEZjnU
bJVJxQ4UcGRI2FZgxiniIr+6TGnItI+wTb9WWEq6gFemAr/+ewlknEw6Zy2qKlCB
fsnUqBZ1vwDca75Kp3sQETwgshdyi7bh8CajlwO+cGX7jX+E2UtSzUmwwBL62RmB
hp6XEupwmnLBkohrIHSBpKdPgKUX5Xe+Jj0bpS48yPOgp/dXb+cVpFyGgdGgneDJ
PHge5+Tr2wA0t8hvvHDCPYnin6VFGBckJjg87chhhXB4AZoVPiucqdNPmqR9WMsk
kgacHFH8Zvl7dcwUKFEaS4w8mL9TtnxTqEBVzkq6mlO/biJAsmR5fmZMRujxmzXw
cL+nhTzXMHH9GriG5NPRu9tkHeZTGPXHmrw+cy2oI9EZCBqU0dCsPh6+QJGJqaoF
10Ck7/r64oZVH903XaAf9YRpSZ8xgrkn5/iZoo8bgO1s1Zy+PlPs/d4M+hRLogOm
o4Mny+eLQbprq2qWqR4Xk3sREkRPmDg/h3WEtUb+lX5oweimSSpIC2i1PY0z+/4t
O7SbxLAFC31wI9Fh53ZDdqTSwwMFYXtjX1iCzB5CG9ckdjPKW6PMJXfBRHHPWANq
AW9PbDome5eH8kbdRjrCLXNj+WYHdGh3qE5TCKpHLmQcQBvynfeTLM/XyNltF2YD
nHY40PkdFcTnjZjeC0gYVCKXahWJ2o24qTJ8qO2zXSoFViztB90B2lrEqBV9MuVH
ggsOM1whcv5bi88/Zxlk+SIcILM2HOOJF+JUU8ovZTmJM/yDUVpWLsyfw2E20UNJ
Ne7H0p3rbaCtMR4LoFkg7Sj3JxJW5X2Wxq0AxHTcOU9i659zfi1mZCGOiItmPBX5
lCBteiyM7lq570/Py6duIswbC+9jiIwqqeneJXKcbvQT64/DdGPhIAkCdOAazzjA
xrVCh5UAqLox2l68TVocvj8vo0E5Y4NIzfDDL/x8aJyVafwKVw7XngE7DN/zUpmq
ZtSNNDvuOdpoPu11eI+s5UAec8Sz7L/ScvQnq1gaqJ59QfVbmo5kW2NmGdKiJIog
R7ZzppNvgRPmHtPuGa/GDv7wxHIcpRF4MFKY30smUJ1He/3qGBvzPsY7/K8L5wMF
S+XrwMUwmQrs8IlMGCmvL1NKA8tLBF5XTR1NRcG8P6G7/AwmU9ntWll4OkwO35OK
7oYzTK2X8K5kiTWkwQbKcKC0vBL3k5jrckrl+t6/SAw8pA6ApHQDyNowco9wqo5W
av1p3h2QwBOtShHT2rInqW34rceHFUXA61cRefSmOw6e3d7+z8Rfk3/Yf9cY6d/c
HfRxnJIhuJkI8GJEXxO8KJxeU3tsM62xaL4dX8t34qdcPVc63t/I3ba5yWqL1OJz
AOA9XeMU8qy9J2iLuH2GkF16g79uR5OEk0mnl5ZVBnFuF4pDSoD+kYbQBILIRhB9
GwlB8ZucSpDFUOBLshcJT9IFs/LB6ULrdnq1W9au/Mo1W3QPi+c4gshQzGpgocd0
D4OZzh+BxrxsOOSNTdBZhn6hZvF3pPOxw4dGswQNUqFio09ltxkcuYpfhaxsHw7A
YAaislLZaj/ai95IKLWwKCEBlNTyssw7HJqHLf+bQsNnU+I9N5n010E9wlpc05ba
C74VK+ZolSpgewY6p/WRAMPwT/2TlxI35QIDjehtUImJoSRLKTnKiE5hMqPB93zQ
C0amwYNQEydkop82hQu7jJetLv9N+Rg5gpS1KY6cMw6GHWLx5XWK2hV844YM7f3b
L1weajPDOMWjLZ2kf5Ao/lhhK0otYuXCTRWfv7EYVUIyw41LdbY/gG6VAXDQPbEU
7cAqhEyWhzFnlioxLnUrUnauy4tQxI+HuE75GZhuZ4vvjVaeAhcNHhopFt/cr6HI
vXQpIdFwWdD5D7YPVceen5sA1Erch6Q1sujkhQi/UKcdie5nnY9GksGtUsceJSco
UPX0cT08FE3ztRDYrVa+AJj7EsvGEOv4ac2GFmJZvV4B2vcmGt2ro6ngo+YS/UiW
MOt8WmDYqWT3/SSQfQxOTKxPBafjV68Jkx4n5O/tVq88e/E075vU1lJy6SJTLoiT
C1WOle5WoRiwzQTDIp2mKOdbSoCBu3mq5xi0V2Z3ewIK0OyIF1iwc8I+QuoClQWQ
Qrgmoa7jJK70g8B2vW2uTROdc8rHzf3VxeYGaHIkcHldwZQWW4OYu9o1ZuLDIYg+
k7+D5xHlMYegcCIJ86BY+8dbNirsirR2ss/GgfFjezGLxOma/9BkEvAgxOgmS5aX
biEoY+LMO/hIFi8Gfwd+n0QdL/lmVKyiZJvhEho2AOy7Zqh3hGqUM9OmBt4nTO1b
WDzPullJSe+2bZXSUwfGp5xZBgjfktBxCE7nZllYLfPR/zGgTyLSiNuC+OzDt8Sn
9V8D+a+PzlXyeQsaxjPuoD8nNuwBw4e67Z5JL780U2pH18wXvONtSvxuHOwNW5aE
BCy4QqSy/NN2aXqNJD/XawWMSFwfuPvaah82Y/fWEwd5gXatQgnv5z9kqFjc5+uL
pXIv9PYw91OxRYls6rm6Kvg7Kf9gyhBUMvE0tMJcRpnTaq4d46YHwd2qA8716WU2
Bdz6CgjE+DYcQSxJ31Ajg1wtyBeZ37iZWsDQ+Im6MXCyhg/iPYsGzALF1hK9EW+J
LrqNdH4dy/9ajMxAHS5TtLC2Stln510rA1ze81gUhkZd9PR46mkXIUyDj5tgtad7
8KsoqDtRF+JomSfm4MJMp98YWwRFK19gakSrdkGYTg6uQNWiYHy495RRYKg/Ga8j
hZCxhLLXcvjC6vaGKDI0Q6ynSIeM9aJlFUuaAdhFnNOej/koZTJyD//dfMm0LyTs
6fZEKNy7dAOU1Advu4nweyCDgjCI8Nfik52/2GSsqrPTL4nKJoYE8AStHyNuss6J
SDOk6DEYfFpLMRqukD4nRkjbTv5kCRu2G78W/Z4e0BQG0TZDsTVHjLN9qK2JobDe
i5DYE8LBt5tkM2NVkAl9TFUQWrT4waFenWxhERd+NZfFCfo1Tz984dKJ4+MlvL3F
OfSCAYw7tfaCc2lSCAUzpb+PsXlAhzrZ0Gjknw1LJRnekrSO0+CnzG8eUstDHLy7
gZIe9P0V4D0bQmhr+HsezDyaMTLP7kFeag0a0l6z1wy/Ry6hj0s1YChHsWwmRKh0
S+w9BIvg7BMUj9y7vN4P7NjQVZABf4UFdUG3XtSsFKLfIzEbj3QwPJzolClsQzD2
RF5UxYLwc2+uunOe3SvyH0DaPprZmgvAvcpQ3x+qYMyPUht7wi9KQM71LA4cbTEH
rdhpdczKKGji/aYlceZdjTmkl8RQOT/ulzKl8OMAQADN+dL/aMjzhqaM1WZCifyA
D/YnJSGz6vF4WdVSmuiXLEQtZZeqEt3OYV53VnXyVwNlpz7Z8aKcsvdlaB2BU7TM
zB68XEoHkmZ6E+1NuFvF5T/a9ewUUuMeuIzHt1/n7/v5ToCwTjhMRBlukMF4CVIh
Rr82UZmQb+4JMkFsu1tuDHFWRvflyeRzl2cJiH6L8169dFfoTN3McA6QUSXbPhou
eAnLVVpRDxjlhoHgkpkzBpSEEY4JsuDVKfEZgVGLhdgiDBMr9nxXuxTrkHzIv9hg
LV2RKHBdNmr1571o12xausotXewR3qDZrp9mMokGqGPo9TQZmWIb5qGmyvyiVdJR
Gx7z2kyDtOD5Q1mrFr1P9vALwEWQvm4zvpvY0irjMe13krnOldGgS80xYo09DrOi
sJp06A5Y39SHwp/UuYItQTVT5TO/C5v/EiXqV8NyDoqkUiI+hHLEM9sB8v5liPSP
rNe88fEb+1g+vVsWAfFZFx5tUuPjwrLGTzbO+X9muEw+IQ8yRvuQMODnqr5w++9d
kB5H1Cclo+OpJ3aAqfc02hLyWVbiI4YZOAa0DlcOdOI1gMwQDPUDQpdiFoEAA3jZ
gufjnJj8YBzCu7r9ZG3fmp7IkO7UvyqMYUbt2o+0axzozHBNJ/xnusL+S6pA4G6f
ZXqjc8ghlLVa8jSZdpo9uXeJM0F7x3r6XCmjn1aQCPckYla2hahZysnGZDCHjhS1
zHudAzvpkZaWD5u6MTLd06VU318te5s78Bo5JeaxIWa5/fIxEkHuZGsc7BqSgoBw
Ps8Gqp3tHGudIR7187dAlbfUhIPOquN+5kECf0YRSNNnwBzd2SbpfMAJtd1EHzzm
UXjPHZtiPJGWHK8QjENopqGwdTXq6WeLo0XrChGikvnjiErkg3lRpoK5xt2Djc7t
k+ZrgqWuwUjlDQsZvXKoWpb/yUGJ0tR/38dujBdkL4hp7ygO0Mi3wvVFHTd26U4h
Ay3eKregjx3/lgttUvti7CXJWDgVNPfq3elYgr3jxxZD1VAJgaMFc4lX+xSDYojU
xEP95jlnjeqGzLLg6lFpy4MIMz4ICHfnvzF0EeKP3pSQ++lUWAO4MpxHy4ZIQzO0
pBBrztOK22I43VxttdjJN6/2PYEPV0aIi1xz6+IfiElVMtFUTGz1RZeQkrgbimUQ
cpyQvs/Kd5y5j065nVcf9xhQuCGGVEOl9CoqQzEBz8t31O/5oLbBHp9/cBUdPmq+
BAe8iBB9SWCaXOqD7FpZUsgiHqxGy4pbBCMzg/rq3p4An3FnsyLkBTuA9M+LlFWD
tJ710FZ7sX/qkH2lcryT1JZ/atZyShwywJSwmmbkQcjhadWlrKPWfr8GymjnBt8z
Ng+GLKsNtAtvoa3xT1DRm95pG5rOq4uwmhULNW3WleFvK81wgEHJx992wx2fdCSk
7OUJt8KGRaZZAY9xeEFhBk6/+MVwcbQhpo54p/RPbsf1aSpkgKyRjkkmPp7C4jAf
jrSKn+FBE5GXG0Z7PBvxFURMI5WLIfxnjrypmmAkTWDVutEOf9RgawV/rASl0b3P
3Gk4Fk2wNCehcP2PRawLvefZKxpkWI+vfBZnrx1IZ8ATddaV/SXxamRkZS35/YyA
u/TtNvTIGU1EBVtD4xKwZo730rT8oQFk5pEbimL2x1ODMiugYGM2M87Z1dcetp/C
4FOeYkb/XFiaeLUkLTraey3ZsDzDOiPOo4luIY+PVtha42HdzeM63ootvdsA6Clk
vawfVlwvSUMP2MEM6aW4iWP0FUicPF+LtjOm5jITq3tWXdtvySx6d7UQSej51PZV
SO5CLKMUPOd7Xu9XEKfuVxAh/Cx2BOiS5MphlBcI7E74LFVoG6AdOSKuH1qU1BF9
Q8sDcLLSL45OzlTlIETfPd0mDRFoEMgo3L3DN/69HFxGhOT1ONndWzISaOVJzLlJ
VGxzHlmM4Za05SodmMY8fG7o54j5vzDso4KoSYOq0EHiq67wqH7Jd4DY6QC6HsWX
WrtFeUvl4HebC28vHGoW1XxwolTqIgOih/dQLsk1mOHqmnVLcFc/jcCUEnmabsYw
ZqmsOf59kQ20CAgJHQ5VONqk3tPF9sRBkuP8aIHleuswvAdXGNU/FivILX1coJhl
tOx6Y59Kr1jWd0aM0jjJOfejqb8JGCC19i4C9qn3dpBNjdBtPys4ZEDDlnJvsoTX
5qosEEQW/XLS9rRRWKE0S7reTClT8v0QuQ1kODO2yXaL82Hn1wL9SJToWtSeH+HA
wqVbh/wGmbhkqu2Dm5d054hnEXAJZbk5s/KnqPfiCQFnJaRODLVqyUULonYiML5i
bnURawkBSlQcbFqhHApHMcX+JMkRJRHWNn/O0jWU4Pzw1CsT+7MdEP2Z+V1bujfB
Sbjl1aRS3FfZ5FJWEBIwHAMeCfbWTM9O48oDCONTUlgDwN6bsdKj7D2UevmrMXI9
T8QnVQyme1zsPZMGLGPHwCrMtkdw8Go8pQ1vUuI/XhAC8QVVP/u0nO/ASUOeUhos
U9cskJbbfH9SIaQK2UZqp5BClNZ7ypFCP+/XrGpzD0suNABmbXmPuCiycgcPEQgH
31zCDsSa9rS/rcS80NbH3wZNUuK/Rn67evE7YYGLeICOIAmkFekIcjYLcSm6eD/7
vqfRvCBHJitK2DGiro6aiW2H7/dp8RP/Us5hxjYLCyemKamg6pSDkKiUrwjOoZqd
8o+a+f7UWBAPJ8gG/lqnEW1Zg0QcpuH9FsTYpnVjRT08bOMV46x6gHagqaPAhcs6
efq3NAMTQCZwziLsLjDbtdrPtZE6kmFDf+RGqoTRq0RD2BWuzfJqx+F+pB5a2Z1W
Ate+BhJE1e1PCNK5QRYGgYM9m/+BcgKOhsWQIQQQqG85QbXOW32xvSwX/LIlGkmV
HFYV6kn5sfBkrGSeg5n7XEGx6hudRRHcss//VS1+CpbW7C43I4/QKLx+bAzGzDgq
0juknWnIIG3iw6j1tDEDCyJ4iZDWJnIL51FC7Ux4saJAYjsZjZpvKHPsZfDmoNk5
ufzs9rjYrsWp//1vPQcnwpR8eJjKJ8L2QCo2JJJIWbvjjAA/T1sBHwlTw07wRZUP
vsVrYXH2cRrY1elPXQKw2Rhbii4wKg/IaU6I4KP0qKRpa6NCZQ4zb0Cq6+bg/2j2
RtcFZ/itACLqfcPDPYxyjj0r90GtcXf5jJ0zKc72te4eY2RIC2iYbayBbj8OcoI6
QQp3apQchLlo/5Yywd2iV9zaeQTXshqxrz/Qm9WKZDswdJOZwqfroBl/bpROm53n
yHjHCbagoceGnq6ClA52U0kM1CR32jaDXha7VzLl1HAvrEFKRir76Vjiu/4PEcA8
lB08IFOwtLy4vlSEfFOcyhkZ3IuQaNhViqgywR7RaKXXf08HYMTes1dZamTddBTb
uzBOduC3pQi5DHcG8w2t7UVJrXAPckEvMMPS2JR9xb4DBbTsWMUwLzL8oCUncIQj
YRIfIa/YSf3XaW2JoCbRgoz72VHWCQehDVADcm8TDe+KzHfErofnfTkSKsg27AC6
TmkxNpJ/B5IswFjAKRzS4w6fUfdmsLVsuF1zWCWDo8Ti9AIqf27xlmd1eZVbDb+6
je30xe7BoiunfVTDqfPSAVvOROo2+bM2fesOgi42X06h3VOWfN2udFpoIZvPn5jD
QWa4vfF3tvN9pUCNlZgF6mGLPzliBGmGZK1gxKBBDR24ibsNdjyqCjrDcFxCS0B2
Smt/Hzpm4D6TiyYjGF1j8cDzIdt6Q+bK1Vw/LYB1iNzAkeelaFlikmfmZ3B3Llc/
X+x5DBPRgYiRYG1ZcblT2RzhcjUAYFjzn3YQuvauhCP7qdyKM5e8ToG3TFUvty9o
rMABJNv5W8+flgUARFy0RDoUzkIvBFXZ+tLWRI4QCwMOuEvFCFBXiUbCW4Gw3gTO
4CxDbC/TN6TlXdTsq3Vt42OJateOj3mMA2/lrMGRcd0C43xwjk5DWkBpu3XPb4P1
w0MDQasPcxVOXJV7S/z3Ev62Ujwl8mvP3FjyKW61lupQY8T44fVWzAEL0Ju11pdx
3hNZoz3/BqSSUwLgQNoysW49gg7OI7m23B4X+uL/bcs6d01vNWWlDIM30Bk7mscm
C6vse2h52/qZJeZN7GvOpfYAc09Tywd7KO8UltWePzF53tyB5KqcDOlck06XQFPd
KqqKEFOmW0DyJpG9rl8STH9u4bHY4qezv10wc77MUyMNmtplzQONC3Wd4ETy4KIA
6V7LeqtFHpNJJDW3yitnvSvtw2slWf3ND04JdADUxOzuMpajflfTKace+xvgz2kR
PPBFYChfF+uom7c4HI/Jcqr8JN5DscqHpgTd3aaIF/e2WeBvYYuwK3nJwDF949XR
J7ISQ4lVoFonqfwwoWQo6bt34KormgjvglZemBgIm2kRsBmnayugHw0H5wL+Hm6r
wJAlH8AbP7uN31Xi3JNQuyXqnu2kcUNqJJ22RRWPodqdrt1iqQBD4xKHH3h8oOSe
GOCofK5Bztc5QK6bXK0RefQAv4HbISY0b8DU/dbG36YHDpiv/WPfZ9BGYcThZTbM
2A+4B9poQxkkAz4F9pLrjLAdUOY3OUjdxVeKjwI64FJPB2IF52+PCUPyCylazXTF
2dyJXQiV1bo7rvC5AEu5Q1ja3+RCmkaeXjzaYarlW6l4DMdWUOGS0A5SdALhhb8G
Fk8I6Pr55IYBC4nDoEVslgckfW0YEJFyTeQbbOvsBpA01NcyPgDw8SN+1GH+5rJD
Aa2leItjmc1JOhgJfydC+c4FG2ATY9ZzoW4ND32bGhRMwRAOGQshyCHvTTmB2oaw
RwZvJSMlrpuhn/G+kWPnb+6nhkfMHSnNho/AaDWgbdItT0OSFrtcjD1sSRRPWnBP
agB6Ocosb0S2akWZFf6Rajp6Ze8CMk3NcENmitUEr2356Gli/QMMggQkKoBEzLI1
dCVmAlnVNzVEFyIJS9qHJLBkpaleEgLbvmWqvGCV3JU1YzlZSmzVh+cj1qW29MEz
/1FFoVqGtNiPE69CTldHC0xDtQqo6uJDQjYRiS+SarEY35WDIoVy4ukQMcV/aQcq
C0HdiDDxlCf8gtVMR8az3B/aOPyAyeh2qsvmcNSHDukbvcwt0yX2jQBI5E8EA9pk
M1gntioOKlQPFjlpNR1ICIYpp4zRrh5/ljGj6/1UhS9auKcgXNt0YR7O4L+LsEFM
6SASRWL/c5pLYcgJGieMIPvXomoKtBrlrEp6ATK4ODKk/ABjckbdo2xH+hAjtBSq
YP1Os1EH6Nu4R/Yx5zxjUTydJ4Zng9yHzPIxrc5rwK/RWtk2rW7P1AzxIr9PZ0mf
WasZgGg7iom+p05qYopm6o2df/RWKpIAR+94ETX6MfGiF4zl3a3j4mJKT1qikbts
sTKl5JV3bhi/XhYm+OTcT7J6w/ykiW6DGJMwJwPHRZexeNy73IYvnXUgMdY8V8Mt
Ub680L5b9tQiUF+9m6V2V1gH2Cs8HBAWD6vI/7mfMCaaHy17z/zZ0pqggmBum48f
LXPeQF8xp8U5y7AbRxWawirVq3fPo+4O0bG7fLfLaZXAPcN/93Uz+kYFmjF8z6/A
vrsfWrSbhd3JsMT3nmu2dXFzICOkckq3svdQQtn0zsVT9tSsOEBo69r9EcB2r+ZG
PNFLtLu2dzu2MEurpfkC0M/15nraVZGw4UJFI5/0yVJqtBOfPa+tP/RqhTI0kwRy
vkC3eK1Ld2FQ7+geZ3TmTiY4zcrXhwMTBLNEDeHCHvKjh1eYquff3kQhvlQVjQCt
OSealcaqwMLWeU+Q1c+y7Q3GGuMlVwTVwwo7UW2Xzn6NOiD+LVc6b96iesbdb/fI
EHURuFOH97ooWywnezuRrSoAvMl89eSKofVTS3pmkuEWnBrHobN5EDfBnJURoFhv
AQfktiUOe4UyeT5YWV5slD3qF5qBpJqQjvhZy8sGHEJZgRhoOJ7Kz5bf5IF/+xXB
7v0v5mGlo+R531YPlM5io/8cz04ERNfV70DVnBOig+q2ZRmx6XGZ2yTwD4nS7yn5
zOaWhvCFq0yG0OcQvfMso+FNX8xYAJ9tKIuhuRs8tu7DWaDZ0EdALqqQVtHM5Pnd
Jrrpzf1+yG1bFIFw6xJYbrpaiMcjqA2rQOHOXE6ntHSn105fxJSnKFzmb3Vw3JH0
ZqdkSbClaqnOqGrgbphUG5455eX1EVRE/nkk84DQkfdIVrXezzxilXzboEO9Ojpf
uqUrpO7z7IZ7a/lCyGt6U8bt4k1iPnQ5Oo7DO13rAiff/qbuwpzDOMWM9Xf1Dn9H
guU+S0YXS4iX66Z1eAjtdZu8srKLrV3x7ZrOChwzdVxtYdAtS2UQeychGJ7oVYjV
Up5kE9l6STXv9b7giXd5XS9yCx7Cs7UhpAmIKx2Q9lWYGLFr4EJV2T3vu2NLHOTw
SrR2CZlRlnSf8mo8YquxAShR0punhv+IFuXDgWZOwbLD9oqMLk7ah974ZfZ633c1
33bXvoc5Tnw/ZCfsuDfbC5ByIViNhKgKoVj+hj7yOn8PaZhHdSkwwkXmey+7G7f+
lBxupMNwcrxcMinAjz9Ti5WCXg9Eo37Dhh0btnzlRcEgE/PE00L6mAczeFSb10wz
xRkl/qwZSxScVSNHe6+d90RvMghwfcXEbd1KeN8jKFuHwm76mLLb+liVBe6GIgVC
sZr21Rb+LYqSTjs3pfqvkFFr4h/EnqbSvFSh9v2SzBY3AROvVD8QZjrjh2BkrsUv
x1BdA3ARoGKc4/HHZsXRveWuVWWW7GsTVVhnowImIitKS1O4znTA/7Z+6FYqwilS
OHfcJ44fcoaSguXIo2MfwG63FqzSHDI2eBXk67RHXFfqEyNniLrP92V+p2YSFXkm
nirnbrntcyyPV8XVwg98P9wtR7GGsw8QHiH1SoztWHIc+jrllrP2sbIWqy9clEhn
F9nKuhJ1m1He5Vtv3lnzk1EwfNBb9WDJu9ShNqo5z3m4xmI+/0qorPgKFTXzqrmL
fjszdRMI9v5Z7ZWSHQF6iDTBitGIP2M7zpK/RCo0skNZSBq1IUKDTWsAMIiji6Ag
WThCbIYo3l4586Hm/6qyeOTTPeDKRYJvq12NnboIvBaeQJtuI38AfnctBlFOGT8M
9xrvU9/gUnJKyZe6xVMpzhzJ9Yhe5IHFp/bmGuOEuzRXWH3TEVxYaxlNIRSEMMle
NNsrDuuJiq29zUQzbGKC1PBUpICrsACdj8JquIMtX3q2ZlUlvvhu4nammWUQBNfU
NKD/HnKhUwuD3hxTZgjjPdEXHkAlboeB1gnttPL2lm+63q8grVqb33e9ZiKAK/+l
tQ1I+oxkupl/TmHSOrrJoUfCvrCWFKuGLWJCLLKkv+s5fNx2aKF5J1D7ue/fOTT1
4HgZR5UecnKMQ/bjO530A6KeEzkCLPmYEquOO5bVBQZujnvVpM4nmtacnOSSossr
2QVTIrGszNVt/ap7YBMeHZ47R9cWLE8mS836yoFn3Oo9bAS++zx64TXs2+jhQlk8
vpROGPJBiyBpVRuj70aXlcu46eeQ8IgjGNt9XwzzaeO3VmH7fZc6EBTy46e+TYv4
L0ojrTWm0hX4/IrKx3FwPEaWMSuva+1xtDe8JO4MxoggvPbr+z3e1iB8to07ATA3
yxm+y1imqx9N6CxXVah1dTR50kW0n7fnaPvEZGTeoBsiFfAweT06rcTZnRjT4Max
1shAJUT3ysvm1f+w1qBw2QgXm5HSr4dTwajirs8B4xo+qes9KoRR4r1tsdlmgoIa
4E959MsdcH1Z9Okct1a6TgK55NC2qUSB7UhATfzsBwaTvdaot/QElq5P7/YeeWDA
ZyvdPaqgrBmY4HsB3K695To+5tEavslg9YqwVcN24kL1l/d5f6zlNLNt6AmmYvKG
cnjIyXoSiU/GdRNFevep0JXyRcnoprB5mBmwfBbUytlV9mcMhsN3ATTDFiJCugjK
cS8XY5dafj7uq2LGcYpnUqbTUa0T7bgWEy9HhnQH+dV6xcE+AJlsnOrhfpJneqWk
if07MBjHaVX/vj+3UMhm97SFsGlpihd3yvomO6wQ3mrpTe6QX+i8sBwJIPsB4YPZ
r4JR3ayzLkOV1syLFsorOanFyZ17DzEDJBSIXY75nsmiaB3do3TxIXkGHrQM1WQS
dVuTHagOy0AwYvCzO9gYMf5UYIb7xX0BukMpiz1ucmffli0Izbv+LgXFmpGzL2I4
55w7oxIxvNg0Aj/qkrb4IcMdJ/iKCvHRjlKp/ZFFiDS0ROY+aC7mI0+Vy9F8m/E6
4nq1vprvcVZS82NfCWUM0qflNcyYYTt3sa4ebFEXP/KVRPzTCCgqE8+Z3pLtfhCj
7q5boiJ/eYzZz+PcnG55r3rVSkjF+KPfqtqKG7g1kNE0SxUDw4Vfu3j2kFydxVw0
82x8QAopjs2888vk9s5VyEmVH3bGkiicqgJBIBcgTXpv9g0nO4dOPMpXyuctze9p
Oe8zZE974H2q8qwPspbiPxBRMU5+AD32+FaO+NDa/VNd6B4SNP853cuwQ3Of35Nb
VIgAl8dOUsxTZKRSYIUW0RN0ejJhKGpahUR7lYE2E8j54DHIkXzrKa3Tlft9ebnc
x9bjEH0Mq7UIDNftLLdg3Bi6e/E2xqbsvxRJCi1MTqxaTnyqktm8zT0Z3jFSiW8W
q9K/TC6dI9kL52pLVFT7VzK04iGc/LkirtlEA7/C4UFqU2EtFpnnK+oQ7Yu/ETDW
g70nY0jSagw9fThz9xh4ULeKxO/JEMVXk6ruW2c0ij4xXqa6F8LRm1zYdYNOC4WM
nwigMWYGbqG7VgfPtnA7IddiiHCtGdYdlxSp9lOqa9/LlbteZxODHKOWiL0IdIgk
Ow0ZnzJlipmdjU90++0FH6ip6USVeM/AFNWio8o8oZ+2wcN1x82mjYy53/CxDnXS
YDLhCN9uoUer6c1sWHNkxSkF0YQx/SGU0tCTBTRYO0osNvHQGH6CDCF38X1EdqQq
aLrekToKSxeoUMsHG2EPsibROL5Orv+7ufB6XPW8UusBsxo4YoGvpt9wyp5p2w9b
oTrCTxBU5z1G+Rui11bvEczFCri3+WZAdSF5Yx4uLDGTzVYQ8IQYkR916ydzjcRl
LlHcgApE8JONNVWBV75C3V0eEUEo7J2mrkUfO44rOYGrAUvCXDmQIg+1C0kS0O6L
nxg8oNBbCKjr2waotaxEiJaJ0Ld8NL5pYuQXCddnwQVKa8D25rpVBEb1OPbpMWWy
PNRMFGHBIlPkSkB78WFP98TKpS4mqsTAK80RtKMBAMbMmr7OsU/cmuPF6CVFQ5Le
MnqICltbquVbrauxNSodFogNRu9P2RH6mF6jsv4FFXcrL5S5segqV1aYovjTvUsL
WWXij/uDotK8qQVcxYNC/JffcDfxfdiTVjAPiuBjDeav62JHYWGXEHvFTVEGrrv6
eofZchNyyNSvREyA4kjOQCbXvm4b/CVz+WI0k3AbM8738CDYk/83wA1E0gXYuzeX
6iMLMMdXUhnmcIcvAk4WRRvAKo128wwIFOmNVin9qslW1GxCto3Yo5bHAwDS5FBu
3f05M2Z1xf75xmJ5GHNjFofeZh06NREXcQMxdO/OEcX9CpY51WXAnY0i+76QnR/l
Z1DJpNMJ7+uzlju5whwrPnWQ7KB7aR0THNHALpSLp29psUKpCAPCl7V1mDBVnrgS
8k/DO8EZAzJXajSbvlNWY40y/jv26UojPHQ039007OAoqIhFATA9TSwwO4ZPRR5Q
7lE2KofdGeckJVTjKOAFYpEZUlutOz8YHJmg4tZANHUZWTmMtTftcJ01nf1K0LNy
HXKBZ1ZaxnyiHB13V4CjoxMM5SjkCth2Fv1y9VFHA4CzJ2MsioiID5LtIwLkqJC7
dQ9obPz6/ReYS9UnnE9yw3tkS9cgsYUSFl2TS77PO+OEVDK/U7rtc63eoIoJjxHl
AYTvYyhzIsvI1MXQW5hYVxZHFtZzKd6uNoa4X6CiQbW3hKu+wWSh6iNy+IV7BoKJ
RHk//FK0orw+hm79A7RLIY/iwuinLZ98DlbxuHh4ch+EFcNkR6tL9bz2j2uVONyn
Re22XsC18U27A5SV0ZmUvsjYqafqvqi9gbb3YmAWV14O7DzdLn5wlxpOHnRkEdYG
4TMll9V+1YZkifgNf33iIpRxDOpkKk/ZLCAKCZhfm3z0iKJjRad9VScpG3+74S8e
V0KToscQK3PpwJuIgxLDmA6sexx8oHMXGeJ1ZQQkj9CYKq2+rn9un3xlJ6Q+Ai62
+h3nc3asRgPSsfqznWcCExcb0Co6XeQbfWg/D9qKbcCKuVbVcWeZCS3r7oAKkjPJ
yP/yL59O946bCIIk0sMwuksDsiRI5vUgZ9ESmiyzsuOh+3/9miA9oxpA2GnVpgfs
rF2cScwKlv0/xbSr2A79RLfH4dzawDQtOWclzTg5FZfL6c7FCkndz4yf2SueTQdR
WbiTzYr5NZDNbCShunzEmGL8LAfmVAioWu3gkbz/WyqdnvJvKLpsg4bCj1fT/uDy
9XEBbGo8AiIGD1Bht1Wmn4F0WbMRqoTsaqtuD85kk2fhHDpOnREItdJME/HL64kT
JIsuvluR/xwiizlIZSw6Y/wGxFbObyUep8GMUaIUf7ZVPWuZOGql8+jTZsuQQmSx
bmqFNlxYQG/tr15c0Ptk1u4Sd3gisxKoCtZzvC65SuDx9V/JioCdcr0Bc7NmLz4s
jz8Yy4tMbWzHNoFtAcVZEofsS2+1CFb5PBg/KBFnUJ48Pc9xVyNjM1nC+3KAtJCY
eoL6PFNflg4nSwUzXZzkc7Q6RROEjyTbePeQTGMBAFwxTVCWcejl88nnqvFUQICa
P1dxQlaQQO2Wjn65sSMAQ1n9RTQaVIHmgcMQdKDrzxOXok36PKNgiswS45jCYIrg
BrMNhi0f+A3bPADzbvmqZnqRKASc/laeYqNVMzZarv1mpjFT/0c5T1YUB30JzU0h
IwOjyBZUfPvSKCfE8VVvpaZi8zlh76fpZ5evPfHzLeqMPvvDtKfH1vhg4Fnz2sO2
9fwdhWCSorW1etj87Ta/IdO2EBjEZug7GuDMDY+DXB4Ix8Qul3ObZYcX0R/I0pV0
tRWg22Len4b7AqVQqe3Oh7qLsmzytH1xJ6IhT7FKL/l+D7JBB18Ny15CiMLvbf/T
8J4TM2Cnf4hTXODVvBlaDSY0feUXSpWiOoUfReDjIyvYnEYzgqscQ4cmGLnMgWk8
NdDToOcEK95jdSlceyJg2du9peRGoTMBKzAcdLzHO2cSGikc3EdWpOzNVQwNm7BA
8EVRoFMogSLSk5hlboo1GASDHLqQTwRKdCFcB1oKSVxmzM0RrwwXTil71aNKH0FI
9HJOm83arkT6X3aqcDK4isCrsEbLXZiGmqDqLBqVeadR7RipTN7D18GZypop9bEi
NNT79MxTR/m9+Cew6baVXBZqqTHA4ZIKBkbdkpcu8IJfP7REOeuZBeiHnEPlBu/G
CMXA5VbuvN29nqpc6K1iE2iCxNkI8KekIzf7ZFiME7oeMSOj0BnvpKTJs7nvU45V
o81RaTJSq/oBjQM8oaUpRK6w4kYKjD2nNZbZkedzDEMXDX77AA1zpoMF5AYXAcz8
FynIAK2zMpegJnIzz9GpC0qjeywz3UN9uMLQlGpElmWqdHcWeSybYfvT8nHQ+EC3
e/vfVzLcrWfWcNzws7Hv47dsxJ38SRsOFHdTHbFBMYGOP/pwSefVzssElx3PBe8M
cZw+MgWrIe5FRECkwec2Fg7DQRwMsCRF93IluPmE+zIbZoMP0q3wsghF+tg+3mg9
kReKOqk8QR/0kBsGLrudmQkKq7Zj7dxYql/GOmqPr+jF7upOMpFk39te5oVcfipS
xoDc7RyAlKIyeqlo6sH4+UNyGEq+5UVXf8uqxv0/73zcjmqiVs8puN99sCJG2dLQ
4EnQBXgc1gGLnlCKGzOwCtnsmMF+Bo4sVgzL8h48PVDoFL1dzY5uYCHogu5gn1G3
8Y1LJh9IWu8ZPEINlqE/qnyzSCHTFvEn2MB7KCL92lvtuqEywNRCSWZL0HVTyQgC
JgkbEoIteBCNpGz2muoTr6Rr0NFrzrsvBlQs/uO4SoVcOuaS65WsCydLhv79R+qy
jF/bg2EZN/y8sMvFFrZTdDq+tc5vL3tZPmljzC83MuJwW4pAGbDhlMuordIkvHQe
tcXZA3OjHkxYOZbUuM534LzD2sax0AC23HlOPKM/0+muURYT+FIR9559V2jTxQYf
HHvxXhqLzqRMnZNEZqcVKUyI6jN9x6jpKgehTXukjKxV1W5gsivNVsFxVfdlsvaj
nO6m6+cfRfLYd8jf0TeZQ233uGgE95Ezw5IkIPR3NcBkzk1spVS9PU9YC9ml7Wy7
SWzVDUnC0NeonfXzziD/DLWTHgy6avtixR89JM8cIfQTnuH2v7gzTLlgnhtNWYbj
p38GS+zevCxmkedaRdrpsmoKYjALmb9r49bB21rEMy0ed0DxLnxv2uOvV8OU1Dtg
fOOa0gN0TdQqiFhmWekW11lXInBsg7LPURu4sn+/R7fVTq6KnnMwdRFLrHHIAh7W
5FLSn31hZpekx3DkzV0vCp3humD0+F1CeSdde3lN3zHhqsRKL9b/JbHOstGXzx8W
h47MBc/sjHA6T4wOdg6kqrs6j/gX0EE1nZ2heY9m9CqZM6hKaT7yChgZvvdB25zJ
5XKSap9FcI13I5KHtwoPacvPbT5jpYKXpCUaZv7wtCoWlpZfLDRV5//+fd1x4jl1
vVIoAWs2XafaStvFxfuutYeF0L35QEMXhm/P7Ic73eZynDjxcgSFb+y63NJZouJZ
RcY/h4jboPuf52502HjBtkYgrthik0GbIZNS/6m5r51ADI0bcZv5CQqP8T1tLJHt
FY88zr3VTr3mJ7XfJrCiBCkVjtjFpFwCfJCa4nX2sl2g9gHiJfyYw0uZ9jDWiDee
8le8qiQZb9sXD+zmhGygvYaJ2q+KjlJK5eiuNWCv98S3Qz3084qOO3gldhn14dx8
EzWE7UW2brAYTtA3n03M3fGkTCWmGH9QnimgIiWOWjKYNCY4eqxn76I0fvmiwCbK
7u0gYTwdXiGH4Xv8t9VaYRdLlUHZy5jpiXi2XHo7YHFM5MZusbSwb9O5oQzJcbl2
cGYwHaW2GzRlB7QAu2bxNlpDtN0AaBDOih2bWbLbdCli8mtbXlQ7BHHtqkd+P4qo
O1azUFPvrSvBJso/1RbpA1OyynrDaCewkDTHnFsB/dUvsY9thi6GBE1thyDt5Jcp
MGcYRFRh3iKkPryczznETp/5sknNgqR8oDKQueI4yeFPoHqY7kpj+ioxOO95zgxo
1Q7nYtX9B8ifFz4bfhgswyTJJvAE8WRUWrwm53mGJSdOhtR8jMmD6QULn9ap3BhM
YvFyd/S3dFroVDFUP3LEjZNcZHVec1KElQtSR1TiQ7okMN0d6+zbbuPwytQqVXsp
3JxOr/yPE19eRwg/2rXtRsU295A/VAPqA2KYzz6gBJqKrjCP4IY1dN5Hgq4zazjF
WpvdCqgIwwSz65JqolXRAaFD8KKFoheyUZWoITWZIAMQK3j/5ux9HQGUmxg8j8Cm
UWpCT8U4CTV0UnC5A1BScYiNIdiGUc+pfctD8vX/0qqx1YgM1E5gZa4Q7UuyY/jw
P9T2ocAM1+qYyjO42gs+0YcCIIJZz3olmi06atJb8xPFq19AWQ/gzPG1lTX5VxfP
1v4LUI6dbgOvqMFOFgDhkpyhD7CmwvRswca8rtIL5xMkmDqfKiqXgyNeRAoyThf1
FyivWlOy9WAsgMsee71hz3iBgA15cjFy3bcUoqU9j9yBl+ZHbnxWbuacLb9yqtaH
yepjS97OSlvcgeb99zprPE/Iqkb+pvjiKFpKzl4lKNfnk/rOetmewKmqh5caHPbd
IEoOCwf8uoFt8SwZhsRIryBDLCutf7wNqPVWXQGJDPAcegn1pqVQgtMEFh6JTy1I
f7pl9bCEwyyn3XPAUq8xBlHJsbIFD0biW1255SvGZnyOlQC/H68XoVib2/nNQ2Vf
/D/uVa2rUedS0d4Yo8Ran0GilZogcsjgv7uo1QNv2Kkm6LjiIZzCUBSe+B6/vZML
KjY78Fd2RFWOMwGO3odERGFO3z9lCANIoFK1bdKwhoQhXodnbqGRbKojcSaSVIIW
ZP4qBu1jVlbcKA3eP1OHtuz3bfqKUG6fCYOsf7EGsCVGvOZM/1X009XgYpMesyqh
2C2YU97tEWZa6wwoTVc5kdmi89vmcbqoXUzOuTBoZB00Y8AiiXb2UQISOfZa+VJA
vmZjPgpj82mWSUIxk5XGUpV8a7kQ1e083+At7fuyuvg3tTmHTXcduMWU+rZfS+nG
+yYYAG77+qb3Y/oc0tcobNjrmp2yoIJQC/vK9Pg30mh9+QqQK0VCp30O1J2a/9ik
1Q2UHkW/JRQr8rFTh+ZNyAat+KJzkR7D+4elENSYfkdq8pSaJy1nVBIWU9WMMblt
sX13cTuREzo1oDg/axQA7Jdvi/tLKsznRTuNB4v4kmyeGeSB79bu0/ULToSXhMFt
BreDcGHv6ORBPWKh3TZLzjN0qcnDhbSFEnGkFS9BxlFeM2uUlfHKJX2RlN8rmMR4
guXyiGKCNp8xG6b4yGKxA6e2IxoWSw9qGa0jpQcW5/gA6GPBi+8+vXRt1VvL+pJE
000rcFeT4WCcq8ztVsUnjWwG/Km2Lf5XEpcGBoyT4BVeQ073Ac++MaK82xoXEhhR
cB43UMhc7V6UA31DASTdErXRN5nB9Pu/v25FWhEFdPI0oAH3iq+XMwK6Eefg0tfe
ZosL1sztP8fHYwQwcpk2aKnUUuSIB0hXAsUKyc6ScAuiunVovLbFU/mTPHdGOy2y
plDt26G/vJR2H+/0eGVpej+WXFOEBoY2O13t8JjaNNAHZSFu9QDF/8jSlqjqsv77
K2oh7z+AwTVYY8ODHHNhzUIUw3qK37rN44ZRrjcRG7456BvOzg5QHtRl13xcpm9L
oJzy4ZGDIkDpiTYZnGp2cd9DeqbCFGxN4Dxrh6E57+cbf5uQCPRe8PFY5xwqvgoS
I++mP066O7cCrksKUJ42eJ+9QxIsm9DoJsSnpLcOkjcLAxfStoPkd/8VOau+3pqm
l657xUnwbcIkL7ixHJDhU7yagiFsLgrFR4PLooMmD43e5cSBa5zQozqpQJI7w8O2
FTtADoJmSaeqI3CSkhjUgsRqgXt7o9kknACbYc4d1opQJdGk1Rjpj3IoRb0wJFB7
MnowOLkTi8mMF6+AM9F/I/3fX34Nc8KTC69y5VNRqoRqXQD68aTdrGaxUP4Z5Rxu
3tJctacYH/z/VuU5k18eAWUuCH7w5r5b7jrDnKdZ4AfQojnEdgBrbyYDv+eR3kCG
Ez7IOmDF6NEPTY2yYKyNk0mj8toDwg0WhrCP5YVSxIvaCfHazZdlEdfvTPggebwb
Cb5/b1TQsIxsCJQPToDWGcQcrW5/yBQTGPoXTN8niM8stDQMXhcrxp2cIvBbCd5z
080y9OsWi1pTZgw9AjyewfHI4EgdiuOiiYrC9AuzKguAUdsji61H0Yv3zsA1G0h9
O9RDckvXI6SsoR2tO7bnJHMxa6QRnXlzPFpP5K9tQbNXlyQ+TK5rkcRxlFy8KDHE
DTG5P4QBLVGkl4y7zZ9pIphIWOfX9YlRRQPp4NOieYQqscEfAtufjl6oqJ7e/R+U
hSKUIwrsODvYV6Ym/pjCuial0nyUqPZ/2PiCB6OSjOE1qAPKMmFyccfjrEoicd95
gwR7TFU7AcBe5dwJlkega1cyaE5eZCvzLBVA318khsO34r69r1IXs6lHJOZZ05w7
6pja3gth1Pe1eyhGrr7hHGnOUSi3uRwghicUY+LK7Bs8X61S1VfMK62ed6/dMcsv
FuLyQ4rRABFBX65t9RPUl1sSJldsLGeVE0aJUy/5FauCxNkjxT0WKpsiJgb3+Qqe
PtYN5Ff7fEOTzHByoftcGyZguvfoleNNCUaSu0JJ18z6J1czUd81OlBI9fuHStI+
0/bLMvfS+d9PUXBVjvvAYNXxUceEux6ueSzUeXx5qvi6O9Up3shRHjW8wsdQisVE
aD51Ryaj6kihBCuHjUAK0/h5bOTxE3ObRTVXJKW+lr+VdGg9Z0NsiOHOS6MyO2kK
5shcewSw6IjuZwtf0Yj5o9fY/CbgHi5qaiSBiMCWrr1TVmzpOek49ng3oayN2s/W
rjpa6vbbrhrHETbuiupkiG8QLvlCOobcZK0QeNYHgl3L5m9/IasriaOKrmdECrX7
6QuOnQBYBo8C4rzElY02IbF6mEjn0lGHvUNZBbBwZuAF9QwgqJd07ZR0sPkZ22qM
GZV+76ksSvttfm3FZ8SbjhactrM8yfsupHnyfzM13GqYrq0EvZr1fpSVclUS0nIh
RJXXPO01O0VQzlaH79755Kl/jPgduOlaothyi5v45S6z86Lr40gMx/mw18rDAY+S
aX3HYcP2zisWIUgh1AroytPn808VEe0grS6mGWX9JE6KK3qLai//NiJxHFp/o4fI
4BVJWbPvoYEk6ox81sJYRNAFvPhkRgDkixlkEzEIafdnEw93ZgOo80trmhsfGIil
Qst43d77U3MmaUWRE4IOxUNmtPWcq2Pt/+ZyBOTMD8qYAVuhjdmnlONzeinTzjmH
0bfoyklOHdAfloqV5+nZQdFxKonyL/GqT4pk0iEKoHiZ8rWjd9vTh6QiPtfWbH0z
1LPHI42202GH4URkjXQzXkfyQQOqkRG3PBO7TwUTTCNwJrv1Jcqm5SOMjQb+kr8Z
sZxnbCZvzQmpro5Yx74vy+Z08a4Bub6Q/cqX/1WlfZKXMDVvgbZIi1+mRg1SdtxA
Avtb2DJc3psJTc4sUn2aaWtTPx7khDFP3AvUyn+qIHWVWHusXymL3WF02JAkjijU
iWFiwWN7LwBG6rdTM4YZMyM3cx1JVBHlViiKWBFzOd8TaB1r+gGObUkSuLvtDaut
iVmNuzJxOjCthqzcA9kdht+OGlPx8pPQYOFmDP1PfyvIcJrfzrhqpd008l4FsFEq
98ArZ8loo+6CzTbyAaeNtwe9gK7SF9qYxqmv2lUQsDsx2ZITVq3W2RPbgp8ABtcc
Itb5iC70ly9OUHludCCX0Zd7apEHFr2LSWLhOyjRbklrEwET1SHqjNkWcrnneqxk
EYy37lGKs9zAhc4h/vpZe3cfDWyi/RMVAKG75DC7v5gzbLouWOX1RCUfi9BTjkiF
y0NWa7sAt2rzUMFuw+FpiOsPAEb2pES+HYl3xiBzuCzAUk9dHeURKChGelgPO+/X
yjdnUDXeBoKZCOzeNnBpKT43Lrap/2MeTXc+gObp6t/WqJ4sCXVdgBd+ooztryow
On94XeVjHZu9jhICgdCIklo1g4rrcX1RCPjbx8NCq5jc28pOugR0TT8cT0MUWbE0
wheSZc6C1BtAg8MgXn2pZ78Ozs0fdfXVEF0evAx6Pm5yKpxpd6poFF7Qk8tTljWA
D+BTFpC8OHZHzOv74ch2znCCHbZgOg9HkYkEsBkBtFrCn/JVi4wXi/AYGyjM/Vvu
lyRkFIQQeDl/jOkn++O3+Y4YBCFiWTkmyylPljfKiLh5IkBco7aP13MJfwLaNpME
1WaulVp4Ikk6quW+QjD7NUhw8O/aQbvXF923ErEujQSTNaqn3F9gd+J50q+R5/zj
T3NFGhBP+F9YCuSn7qgOUzHQlU1ylheTUWJE5afk723wWhd6gy76U0kGxuHWNlbN
xAzppWBpZW8FPWrxdrPH4Ghv2TJO+z6oie0ZkEXl3r4RXgFmD4j+MDBsdBoiAeGD
Mgi8CKjDumQ3/RlEqO03ugFJgWW+UP4qKAoOB/7cyVQYehA60rjsoumaOpSAkTzh
VKM0nuhF/vPjnbGx1OznPN5GzOVVED1gu5YLWndPUhxNRIg3k1NR5hOgSh1hjhGN
uoeCZh7AODKa6xKZbEZCOz0Pwv651IRpPobhahs8xfIeHE7Z1K/nN1QiHn+C975B
cMEH2aaFjeUU83DdOY3R2iGYTlk2vf/BL5Sq+1RrkeD8aEA7h+3rOUiOHY6flRbt
6Kjx1iwnWCyyFP7PaJ/FWVqPD5c2nYYfgQ5NnHIRePnGJA0h9MeOjmU98+848f10
T1XWbP7f8lSYTqiwBRnbOXpwNLdxcOdMlBt39zdr4c7PFbENCJUHMcpNwhjRdUH8
YkuIklKUjdVKoZP9xOADYrWofqVn8CNdyCpZ8hHI63CMgkk+vVLu5IBgRT1/5v4C
NR6KTX5QiklP+7CmxTKkhXvRQNgl0Wg99UW1SWKCPM5YeWa7F+9EjC2uLDm8s4fB
+T1NER6694eSeWVmN3gPnpgtfYEdJ86vGcwxSs06Vzxm2+2KcoGtWTe+2zV94CG9
WWE6n7/jbC7ZqQQSGjYV3CnNKxYefQzALykXts4Z+NXFuGz4KN6bvWPCehMpI09T
nr80aFGaRCG99Ww1vbmk5tgiFui9wallr+gSBLpeN7Tsir6ThNxduwz6xand+GJ9
BbFk24hJ+3DEa9K/cR8VRRA89fWdvyYTem7tknbqyPYpMT0JxcJ7xBVLDDjc7cJr
/PQtxZiFRC46/fxqaQFH3je0BRgvj0UIqSj7+lFrihYaGe69tK09hk4PaEiqM+Nw
QOWPaJMEtWzEtP5eJ27/FIYVkxTFZW9HgnF3XJ93BjG9C0gYIBevhF5ExokluOfg
iV1PVoU1KuW8zKbYm+lSNWGcWKwK35HjJIUPrNiiTxkawUVs7Vua9GyIBlVBimsQ
08PybEbve1XvDyYxc5wXc7mHrEFh1yZmUPxu/22Ddl7y9WS84YMC7TNsHoPDLGSQ
8RxrhwyYJS2pa35S1FGOVFSKPOcI2v6bkXH53YAfMKn8My6wZaPtqRv9Uy100SqP
xwnioXstx8PlksF/iAzhLQqv/a1QI8EngRTOph4gJ/5gUTaUuvvpqiaAVigL+pYE
9UQJ4/qctQyLghrUBN+/c/GyLuHFzKemdUX/tQqTgYDYsQQtsDejdMGUW3I4Mu2i
2HRtuqvi1d5ZVMwR4UVkh4my0qWxOBzfwQ9B2iv2EfduHlEwl4yDFaPpgk4AdolI
gfqfGTdfMSECJ+S3tVTID3PvvG309wF82DmYlmYAHdQNU1d3ocSzDGm+IBq18Zuw
fdgH7VZhP2uchgLSKOstG1bHLYSmOBDWAgVKwTO45J4nsmsBVAPBpzIXUpIImHu9
sHxrloHk3ERViG8aQBIkeOUT026/AuQ2d8XJB8mqd+DY2sSvDBnPzy3h8NLSV7qN
yzuGedTadQjLOmjP6w38I4y375ZGdqZGe4UdpOLIi5MwqBg6xrmDV+wAEI+OCQI+
cjOu/F4e9ONS+g+WZfezIe8rCHTeyeelmOpp4wJgG1cXGRYUVGXTYpddvNvxOZYM
FjtVxbok7N4ZKpN9SKKujMloMNJBNYDwrB0JiAodPpLx7j/sRDz1pjpCD7AiBZix
FS84MQ7A3N1X8YAY2kOD9LFORtKE5c+o3AyValEqHKbPGOy/FsWJdGbLL6YAVAOs
cbuLlui8f3L7zPxBvbI7/z4shwU8YNuuR8ejBn3E2G1R9vVDIB/db8+b2U88gcFJ
673oYKGcJO6qCySCaf09YJsATaNdoDyVWicfl2vKLRfHA8o0EhP8edFD0+sgaH+9
Gztteg7eR0PUNAH1gex3kae7vVxfu+WC0emZztYM4laWcQ/H3pll+AlfBZ75STZz
rnlOGVvpkc/5J+TvdQpk39QWY6RafZeI1zTgJs7JWZIKXIAJFAYJhghZwPz+TyrU
zq6ql6iGfkfHBP/fj7zgWUi/WVpb8Xqy7rVbIL5eK46YAyk5rGk1hoBjLawzKpPZ
MXtXNJw4XwvaR/pXys139Np39ncmF3aiDy42xm9SWdd7Ggn3SkVU/OpAK0Vsy+aK
Sd/1Gdschmqo9xT5yTlbzMpb6dd9kkdaER8r6n/6mSwhF1Yb/RfK3+oDnPzFUB47
Sc7Yb/yAat9Jv5u+0+gnmwqualwB+BI6X2f/+MInfKjqsqxDsDJRh9RMDNv4fkM8
/6Zmw7JSgxyFtgyjS55dtCjqe4/g2bTpzy86DywL6ruh7ZnNEz5uThmlwjdfelfJ
EcZP+plWwBXYxiVEhP1NcsSm1/BR7HPQDJ/GJwkV3M1CJA2iY0nT7OnLe/ZoLJZj
X0pcjInw1WDUv9TgF7ZY6Rp/khsj/xqKzns8N5wIXtRRuAHJKu8JDVJhNyFFK5C2
0osnZ2eiSn0iasJIyLDLVayA1qHyXAcA3ltv8FGGkjgMho/dxUxgxoLcBcNaYVPx
yiQImpiODwaA8GD2KnIz3arfOaBMJ7zjG/SPM2gikaCFWmvpgo6JGTh3SbRj59wS
MD8IMAJ1nOLwh6D9jcgO4HtYW1ctjU8ky0qFd9Nd1bwy3oCzOI5cdt5LjERnpyl5
Vo3xk4fN5LqphTEwK3F3IGdrjbiXyaH7+AbkOBvRdnqDPUXiAF+gg/NGMSfdxm6N
0ZH9DDkbGU3ZKxiTe5TvbTEQmfuurSAC3mpND8rF6/c4Yf9v15wAJT7v6LH/o8LP
dh3qph0zKYVbZQYCerCPFhhPP87nppSMCukJ1iBdEwzazJ1p3qS/j2xaC2tC1sxd
bcF5SpdlZBKy3UaQDZNyvDm9gzEaSXhMmW/TKmUkw/2WfgdAFmmu9SlWE2iReNkr
JJR7pMejUtPyoZLihnY5G6i5QV97t1YOg7VurazTFhHlVav4810pOw8k0Eh3HZjs
Y/cngJtOYJhyeebUzFgd4aD+Oe5sCLVWPMPJ8as9EYBdTH8i8SO5ZeYI8UL6ACod
MYzwNj0S3YWXzgv6fKdrDvxCgwkcZUKo8FmfDM2IHJT/Bl3kjN0iTv/pyDMpkpxO
FB+3nrtRvE+ydT+yVqwP+a+f8gWFvsUUxu7jvT/6vMBjF//yippn8GzSnRhjpBdv
a/fEXvKVF44ElBY9lwLXg5eInbAbd99Evuqi92PAWCoOKOSAMiyN1gVp+CZLgbO4
LLVb4u0OCZNJFv/qVZ/koQG40lJC29LLhX2f2wKfiFOkf+EaaUuJvko66A1TqTaK
FYYDaXoT5J2XVs23KnPGNxKEj+DZZZCHK6fNyAEzOkO6NajneZGtJp4I6Yp26fUc
aQ6DUDabLJqCQjOSkkjlIBKTXtJVjMWky75raMD5Z2eIr+jTACmhuzF4gytQG7G6
HR1rUvVPWLdunGQ3dDhl2rEpz6sqLQbDiqRjDYRBVZyDhklR+NwwHqlLK+0/eMPm
6OuXcb77J6WOuI22jbXX3kOaO5u2au7dL2xoNZdb9BaaTR8yg928cE3OJD8Hqi0P
y/23hvOeoxud73JgfcFntVA+1elylTjEcUyrSNJeIUJh8QlMLWQ5rqfiseksQJ+L
K1nIKekOHlpJ+nE5vCPCvdcV0PutusnNf8DOrg1KWDYnzb2W/WQcKckZAPB40CzK
sRbDAm5OLkHmlQ3gaHPpNulRbi5FDYMaTEva8qTbMqHfIZTvrbFIWPIiw6AzsYHb
6uMW06JtLCYD3YLTj2t/7+bBtzZct3g7sP/tL3TB88I//kWl78p1Cu4Nv4PwKmc1
rLUSGitYGSKB4eKCQuOXMTkaV69hiRmSI0hvW7GRAYkijkuN25tt0mzvrB/hy7o2
VLBqSlKTnEb7oDnGuHyKb1Q8rhoGHIDs5bDfB8rbafUJbc9mpV32S/YxLxTPoQAW
VAvxgdxExquqwWFFxFOk0pPTWhls+0cepQXvXe6T2dpOkswzW9AzeiUcOrrhIi//
ydAMf8tqYJnxYUbkPNeJJaDQMEhi1ZryTXe19rNmjkFGXNufdl+F7OuNO/fIPnGy
erP55DvBQ9ZF8ULv7hGeCld5JJnHOEbrRYi2DjVgUm6APqGRfAh8eMjkpiPAXT/z
GaAmauMA68Wibmz7tAyNiMa+MgdJglyD1wMY0UUfizWphlTxhIMxTX6J5JDjdDnP
cG5HW6ooVEh8o2bHaRtRz0ts1ED1LsVebYtmvzZeKFK9+ab7UaDpp3GhVgjk74Wv
U2e3WrbUxu/S4QMIPGHEF8nEuvCxShraF/b/u0egCs+QCoUBt96O86HKkLBgrGS2
zGnL9mGzWxvovaPW5ispUSu0fFuiT7FyDl1fQKZrC3q64kv6kMudRhmSfw+z3Qlu
A/bQ6EVw1I0b2y/zhhPZONm8NG4NmXs3YC3/u1eeLlUpQSuWPynVStrOK5Xepq2I
GpD37uDND3LQdlrauOAQz2H8pO96O/RKnb8zAomMeCBRRUZbpmZ1DUyRrttwE+eq
tQIa7zsKWrUVBDdT4M2kWDTiIhn2bG124Nznamp33tTtYKhvLci0ScHZdQwd+IAP
qVqKrv+ucR58EBWx8EFv+n9oyhjqWHwEpofUys+sv3LTIrI7elMVYEVYxAJ6vuZI
2qERJMAeJkauSvQx9VoLuy42b0a0H7PrB1rSm9hE87SUvGBLE+o0l4QPKqUL0Hb0
ZwI63z1T9XscltYIeJ/YpQWOaxV8/2UH9dCx+UifLcdccZQ9ercXYaD14M+cWpQi
1iB35CzDmfym+o2esLQP5HBQngBCHtpB8eN0kJfwsFtwMEBVuE9HlDvqZR4vNcVf
FfWcPddAArQVyhjomkG6/LRtR9Nqw3B90Dlrw3pjUPD0ByjDSZhVg5m7esuKpoyO
0MUFc6lKN/J7/RIE091PhlfqVeqwijpdWlWs96GqThG5x/COvq7yBX0hvVyb3myc
3ztpZZqbpWNrkCq0vb/ZUynNycMVf4GxPTAUZpt1R8kqvHL+u6thLn8b4WSEgk/2
g6Xfla0cVlZPvrwTJfJuO6Jkg0vra6xZ0QES9BS4Nk41Ljx7fXPHnPRomUlBWaGV
2DKbsS4qCGeuuZadq8DDl8/HzCQ9k31Cyqbm5R9ZPpGbQQGKFwxxs9X1qUFGJroY
2KJ8FL5Vg+Ki0qL2xzXhTYgHDoZJbC0unyPJGZP5pZ3X1JGCiHrkga63Vnr85RiF
6A+/uXXTWPpuBYE5lMb5zHyjznzOG+s7JX7rfYfls2OiZE/yVxI5ydc8Y6OEcmUk
KdIU4mlFrl59IcqKhE0jAX1m+vhLM5f5kfeTHvwDnCha2psr/w6d1FCUn39yFrFB
jMqaP7jORqsiDg6ihBbIOC6BVGHr7zOO//7CyI5mzaIzLPU3Az3rchmZiy3e2N9A
yA3QWi4HjISu5K2c2qal1x2Bz4N0KCJC81UE++LyK9kzeuuQNlI4RKxUt9Ui3P6V
lXO2GrUI3+ftu7dU1k8rPM0xGNuS4IzyoJ9ovwhJNGVJtV9k8GgLu7hBlDN2PdpD
GVEWyOW2zOBYSG7UVIjXDFh9FTY0GppECeMsVwDgkefqEcimKz4Gu9egP2tcEdVT
TJc5i9V/2VBPCk8Fnqb13PtzMwED9Ks9twY83iJzu6pue8zpY1oXduLH3gyubjY0
7/B5PW4fBF2Rro8DawCAixJBKNVTg33RG/rnrsLPQ8BPv1QBp5fKyYdUN3W09WGL
iIBg9hw0xMbaubk1lVo7e7wRMMXaIMXehv/ssJ8Qn44DDDZFVlNRzcjS6fUSxBeh
o3kkgffY8c/ypiIWaOaUQSVrj9ZXasgkonQy9XuKkoLsWBzPIDqYCoyNNHR56YxB
6bG392a7fkS7NvQySgeYEXsdNHkr1Yx7n8AQYuVh5PJ0HuixUDWPHmf3hAhNs1TZ
VijeWvXuB16w3pUYK5FDJvCDjxZWmuVaK/efzcmuElB38gmQplBt0wLwu0YVjYiu
VM0lwcqe9jqFgl8RtqDO2pFFJKQq49HrCfkalHqpm8azzKxz5YNssmWjPdnyCZpz
+ZBfGJECZvHvGG9fOKLqOQeaI5qZR2rA8INTLFn1nMrHS03g4GpkxKhNXbtBmvzZ
PiL/5BftTlN/Zt58ITS7gvtHg8rcqaaQxEmzKwRd+P2SESOH58sRNFDsG51VCv+Y
pFiMgsAX8L+fdhvBIziJPFuBVGHQK3M1svKh6F4Pu4bxhpsf4eI+pjOfD6GAQKRt
xVogmI9v5yiMD+gV3FxUay12EYM0nN2jMuG906GctmX5BefAl0tjNo0XEf2eIrdh
gQhKvHVyoZ9Cd7e7jbDGCMlfwpTiBiD/jgtB8BILvN1IdVz2PGWUIuo/vxCipiPQ
WcdZX7ynlfAF0xzurZ9UKwwVMM4m1i60F0Z/zpMT2mgzMD6+YXXGxfVJhGsGwQih
MWGfavHFkvUeOBqw+dwGQ3o2eOGAc87eBH+xKLOs5hIxmbbhz1OFlEfPNoSZGaJ8
ANC+AkOVfxCX6thRDa6qvj+rKs/nfZccSd4Lke6jWisg4SQJLmidfMbDEauGRHoy
IeIt1AlQYDl2HhukRa1dgt6WKzhrp55BMEpB2TH9rRZh0IH+8MsSIHFrV6EO7+hy
g/PA3qEHoG0cGH7XTa0+rXyEDHa1DXkz8ey1hUHgayB9pQCRqwrKSKdipb4KE12k
pYQGbX2SGg5Ig7EWiI1VMh/qMvghTfLlP6g71/XVYgG1slGvSbxRSCjxKr7kRkgz
ALd9RCqTFiQ3G1tDh+gUAo0dZrSl4cx/EPhHsqiQDnD8kQPtysAjx2wwE0pR2uyS
ffHUIix2M5FKGomvedWoTxEZ24nrhLXZR8nO8UptOL3t3AzKr8RbK35+C54e0hD6
1FlkdXRx1jT5T1bI5mkFfk1wrrzIl7yGTHHF3lOxqF3q0qZmn7qsZJjs3p53IHOv
6/adbdMIF5FVWltQvR6Bgv0TVn3w8qvhzKPXxxesA1/kYmt0x5e/IzS1VjGzwEtE
SZsIMWjX/vDO/ei88rpdMjbRLlUEDo71U3fk/Ow7+PNI6GGMPYFQJqheC5WTwn7i
5HjOv7MSyyWgZMirfcPSYeI7As4aLDlb3S3o07TpnTNq6JjGZdslQC/K0dGkPuny
+l7W714CS9Fui5JPegwvat378oIqPaW/HzNF3TEFYGAG5JxPkAhdKuzGwwwJ6sj+
Vlv/d3i0m46ARzY3q5xq1bXLVGC94LNPo7tdIAZR+LdPOOSzdH1Om1Qz1I/mb046
mBwq5UpiuK8JE8wlDotWPCkYfBIbV4p0hjT17Yd2pkvqv/ObhKTlJEYIRtBa09wy
claPJvrupe56cl2zukJoXAQikYCpobYavG6SQkyD6pPLZ3RA19hvEOk5bJou6Al2
yXT4v78e9FPwi6X3cGWLbsidgEJAWlDOWHk27AEI1KIzYoff/EEkWlFUQxldKdAt
e9uIIgyNQTsQgLMFaK09B8Oay64srVbtuU1YwbHTAC7TYhHQxPD81h4LG7UsmRn/
DiTtu+P41t52wq5a9dYibTTZhWT4dErpn8ptL0FC3KT3wQMbWC5P6Cc5qICghonv
FHXjGsYkKBo3mjyAQL7gW0LcoBZ4rJkovvYMSpxZhdJBuGNwk8NXLKgOmFfEHFuw
58ApNgcwvjH285QgRhqZ/BpdXxQO+qLR7MdfK4GOxcAZj8t2exaaDB62xQdXO04/
BkyUxE787m1HnWEps+RdACdKKc8LmNpcfy8VlcjKAAcabKfb1rI9MiiB2ywvs9J/
uIGdTTCeDDQR9E7GiYmRRg4PNHq0zWjEv8dEWv/YPlZBm6CTQqleI9GlT8sqEj0y
5rQ1ui155itKU+jdzcTtDmaBFIxUAUafExgF7TKDk0mOersQ0CIM30gds2X6eGGk
jxf3JXMvHvvTrsVaBMG3CTayyV0OIZxFhwlu54pBqblM8kp8wcsiGgSR2CPgsu55
LuV37n7YP73Y0KyTWh/5UG4pIgE08T8ej/USUP5iEBQEfm5xMJlEhfAupsZhgEiY
HcD9vkoRpcoswreNnLJxA8LlhCAkZGBFQfLuVqs0DvVxQ4YroaAI9jX9dcAlJ8ma
yeu/eIO/I73N4RCl1XMnw0mfZbIv36HgIaol28P+Y02pSsguLonsze4+Bon+QUgv
xOt09nPv4cRSvsz5BqG/l+0mYVQch2pnavQAd1EkJkq4FSSTVSMJYqy0ROWFm+Xc
HoqOt7Ne9nUtYXyRRI7LRIExObQ6lQ8ueJ7gnSofhI4y2Dx8N0L1/3l9aFyBbdHv
0aKAJxTIpRREUFa0oQ2DZwc7/lEf2yDTf5XbATgkIqV/NjO7w71rmb5BEpJUa4GZ
ogp1dv4sqcGVh7CPMwaTrx67pzvDP+OUkW5woyAsOQSthbYbhrSP0lyVuKGdT0JO
eBAgiIDS1LoaY+3Vi9Jy109Ap+9dC7Tn9hUGt8aq2DwuUfetAT2vlSc621oE13QY
HtvMr9m/YEQ0bJOzf5JAeHmCDTQ4/eu0622yfhrbpdLlBfGvfGgyHhkboFAXOi5z
RfFu/WB7EMIXOHTHbpo7/I5JObDMqi6HaB/6xzbyQPejnpFscODWeLBvWYlvuJ/c
LbTE89qnvh5cQ4mze7LpsmSxNYP8QyQ76GrNRQcX0DvIOCUa3VemOU8i1HdKIP+w
iEMP+rkx2QFTxHZM0UDJdUtFL/FJ4UwI6st9QfVlnR4zNbTEfmf43KSSs9X9hcAr
PT94QvJ18a6R1ZtMkje4ZgUWvCdJQ50vFyu8swEaBYzIT7L0DWbzQYILoTLEptLe
MSH1UcC7j9fQmauasotVD+LfmxcTW7ElAqwhNCjv3qJTA/R1qLVRLJKrg7W2hP11
ZYd5NUsabvi462ls4GPD9CRGCmSu0DjWGiXlO0WyV7EGb4hLYaWV4B7VN75CmvHk
aaQNvGq435K+0PI5TE48EjgtcInzfxv2+fI0yIW6qubIzfxK+0UXggc+5LbPDmm4
YFsCqkxZwgAPZUP5c1nRhWh/si6gTtuzjddBU58DhiQB3+X/FUhx0IImYZAqStVR
BgNM6Z4D9bqCW568TWBfGmDZIjPGpNTzJh46JrLOodJq5McDWEE4RFlNppeIxxuz
htNw0kxkPggcHZVC+oV7CO7JJNrA/nS8a97TmO2yuakhHLQYL6oUK1hUL2Gsemh8
yGCLltJzHgH/XcZjg7xtijCN790i0pUsWDogynaUO5TS/+MCbsPxEed8eaj+XBCT
QAknGFuLpRJYnb4GfUvMlnpMGY0jPpVfZrsrTyzDRCyA8UVBwuF7e5Jv+9GNztgX
VTwNiLCjzuz8+kxWBqEIfV52izKDu4hU8evfrhZnFSNWhHr56f2P95L+q8ouyoUT
6E+TxqNJD+cTUZeSbaoYxqMLEkdh1BSwHQSuwgf4X7Z42NkN+lx4zgOqRUQbMMIH
HBm63CPQVsfQaH1U6oYUf2Ze+RE7LDW0GyTY7Vh/iMEOn9lLTH8fx/dbcpzAzkKs
jl+d/viSqfGIWHDwEAwExCc/4L2OrP5cWN4CgpX3wf4sIlBG/8UTzVjpVzIP+iE2
oCSnGqmVSbTfA4UFcNDRetu6vogTuj0wwR06aGGllDdrD431+NwOsB9+G3MscbnL
vHifDVLSAuBR7QtNAb5JRR4KHXsaCRaCAvuy1083OVQXmMlZfNY8zYHZSlJGGfF6
WAxhe3OufT9jf7xldlDVwLjB+hKUfYUOMZBkw6CocaPkSsbqPGvOPwn+u5A/rvms
DoCc0bk5CFXoH90r+jgVEdRM6cQkcCwCQkAJin3xgdv1mkx+rFpf2Tlq3xx1mUL5
pBGTEA7ZVpRoYBHlUVvCvEOOwEuwbu//gvpGcTSN2MSpan5Rqzr/oDg7vtY/cspy
VAw7+I5g09FhcdJ9gsFwL7EO5hl8KqR7AbEcAcwBXKm1I6coeTVG0yMrxQKH3bXN
/pCiE6OQACTODArm7ATTnOsYkWwDC4OT7ejnuvveT8NJ9L2CaBOTeh0ITP4EnPS3
LuUCt6KOwNATLBjSc9vG2QmT9hDUCK2hGt6fAPS/rCWTTQ/9s2lqdjHeTQ8AU4H/
O+8LLg83j+RyRWzVju+d3yRUxHljIqnA7lXlPWs2HC4qW0+NCt4kyRevW1wvL4ad
p7MG/XzEJ0LEXxQY4B6awv0kGa3JhM6ysmtB4MD/P/gNcKMCIcHO/itR3/HqwcLT
Qx7NT10V86GFRnN5LTxZ+g7GX/gjhzxwg1VzTPu2lyEJdBaATMN9Jx5hBFMxwwEZ
RoN9xyG8ftaEdMzsejneNmZBRrFZla7YT+T91RVtnuvvEnNJoPBomKNHi2xZnLjU
iEZNTqBRnBVcl6LTbhSjKYnTbLMXvQ8qeiT8o9twTTj1gClRP4EyK0N/PkUwg6vG
Re39p/bqbtKNl/u4gVFLP33TceluzZ+YOTt5D+UVux3AfRT6fLMKPfG7AMEDa7QR
nRgONFssMJqVrpg0gZ2RHkWClqe1brDzFGz1xSMkd61hG2BLQr8H/XXh/Qgf3Xpi
Vj0F7EBj1+P5f7UUV5a1z0RkgjsgJiVx1sNTgTV9e6Es/XIczcX7WWthm+dzBmjs
3vz+qH6mws5M+ACAEfgRWU1gICrfC7OZnsLHAEx1WkA3A0ddCrSsjop30u4Kk87r
SXhg1qG4iRG4wp7ZoZyOJztuPFwy8qJECWm/lteW0iWBmhEZ1ZMjPeSXs4pJtcTO
I7rd81l0YdJK29hw+S3i/tETPc94y4/o9Dah5yTgMtvDIyUOXrP3cJRdKC16+svg
iA2CQIxDqlqKPUNO6/Dyg6+u7rpqzl6Nk22Jhx+tPlGSebq7oCz+2MIJL705jQ8j
QRbh/N5ICXI+WoYm521tXisRC2/WFxfArrKl8qcVg5r0O5dcDM8mZo9fMXEKYBBG
63xRFRy5xDXVqRDt/zYfvcN9PmKiTPxeqQzzxGlx+45IOLSbKWuW4hOQhJnXccXP
13DPmCIVLQx+sEfCwbeliImTt5yLtHIR7i3UtJuJKiEf4gazVBdZflyI5t92l+w5
O17J1Q5uTgiXHdfhiEAwHzcoOU8eBeql0FW2D2zoY3PITXzdTblq2/x8yNhQaYcV
mceo7cm1GCWQnpbcNjtzbAZOGWVVpklU/gdEiASeAyBPhfLnbx6m8xaSgLtucD1o
4nNLqqr2nooVavcNred4n1j6CoC4eanniLrria1DXelJxcC1wOBVyts9kVB+xAIG
jPFmtbfWnBDU5Fx3by25i7VVggcV9JR5w4XfFy2F5g3l6PXXfAXaKgH/HWAJE9fc
j2e6RkLWUCyWDB77l4aDkvFO09RjHmJaNVZo/1MIrdy/gpJJEGre7kDNNIZTiQ0h
L5S6l8jolXBhAuEWOTftKg+suj0vBZhxHB5ndz91lZHitLJVGUCVMLe7Qdfx0hDM
cAW6kqQgrSuYmiObkpR1GsiB8ubBnH9M6W68NxuKSJ5yE96duBZgOkCzM8bXHNzS
Ehc2gaD8zE8MocmgIMwn1//Knw7tLbceYl6U+XQtA/pd4RF33ESHSen0BLk75E5T
LDtK4CAt90WoRjXbrgmKInKJgOvw0Nzfsv1+7bx26HdNLowDio0neDaUyupGx6OH
6EY51oT0lLEObthXQ6eKyjIE9v7hDKUj7nV9eHn0BOsSCbybsMbw4PDb2ZmvWne7
NkakQo77VHAmn+4xgOztBo+5otSmX+mgk6JQwt83/6nC3dp/6z4y3CVuE/7kRbyb
04atA91OyDS8nOveeoRBBfZIFOCXIjEVUGPsKie5LtXkMC1ygmyctNitww+j5V8l
B4iNTZzGtPEmelXQ5/ZwszivMWuL3LcInI3QX5tbWMN6L7wTJ5Ply7xf1zc4WUzQ
jf0bWFHPNQuiK+4SJZuOE9hPDINbpI6WYcqswdSX2MlNouqC5J6BmUG3AJEyiGbe
tDEvbMNAv/LhBYe/keRBV4KkMPBY04Wl4j4bbdUmMg3TVnr9CtogM4AApkplUYz4
6ILGU2pKeezzvYS0nwfyH/PqYOUquAYCQXuoVuV+O/hVFinZzqeVy3PVsrcEvs/f
DevKF/vaEFS/TYwzN8gBnVKEkIiQtenD+9nBk5VcJeuGxOk1qGNmZaSHAu2KmNU3
kbM/gbA8kdkg7/oCRcwx2otMDO0xb3l32ejAS6AZEXpXTOKnZjiRHaNXSP2R3SJ+
oA9WP8YcJPQS5zsDT+LqQ1civWPgO7CeY5E7Ag+FegjM08UjVXrREWzUkhAqqQ35
kD0UrPhrDaGfiksccGrsPpz2F5kFwFMIYxRXW4GV0QwRLglK3/DWY4oSUQG1yLV5
UxGj3KuFWdircBfNeE1zho58gFkyJGqLFRswBmDXb24xGWZQ6wyXFaHCW8w3ZkQX
05KphZJAmP5o0BWgJZVXfToPqYXVrdvuE8eQ4QzMJ51szVcITNXw8tfg+4G12tYi
/O9ciUWlj44ELh0lK2qimOuOjj8jwre+BHdV2f+R0Y8cDOT4kGaf6mq8CCwMHlhm
DW7DVKaKdZLroQxYQPModxs1NEIi1oB9w/IZOVlc8Rx/hEKsy0Sbo6OiSxh/oE4r
8/bb4r9xY1P0VwuqvAsDm0+yruQtaE/mJgi7lKxYZZr7l/8HQZlHtcUxisbFTL54
3+gA2QoVRDeg14fUmubXoqsG1VLT3Ez4iercEQzQdIu7BT66d8LsT3umH9y7Mi5v
DY2tD3o+h7YFU5APz6o1F2qvse6deX4aqxBEdSvbjsRk963HWN6SWe01YeyMmqIW
DGLnxPeAkJwjgGBI9HqiDGeeYzmgJmK0warBunKpZCuPLrH6lsreVWumU0wz+BAS
JtHKTZcwPk3Sl8bBh3KvFxrXKukdTg8j2vSr61qRqSNiJsE6tUly+yGiP36YOczk
TAbCIvfss7EGqGMjDGX9FP54Ttl/ACHTjSaWEhS5m6qauopoRVk6QEhbo8gq3CMo
+uXBXYrzadrVaP6U7FfbDVqN2ORBRdMWXqAsuNJ7uM6yUpQv32cfdRNFB4FxwOwb
eBFcmfpfKui3quDbut0dCydBnnt5oeb9jq3Uk5v6tHLZGMNvGwRa8f94+eU0W4Px
rWHbDnZk39VXBL4gRXrH3qaJJOzjNrEs5yZqP93eoGj9JgEU0b4oZRIycxt9ozSF
OBoAxg9bcQjErr9GIp3HmOBC2wB0K26vUFg8lsHhE2oo9iD1mTVYLfBdgZPBzdLP
9LELJqMWFYG/NZQjsMod0grPljZB2QTCO017fP/jCcS436TvuFuDDkjL4ccVFxdf
AV1fYFxMFHPlJEoknpxjHyr+CPjlJbUxEkJxR/MEVtqWuzGbO22JammFFC0c3jrn
KoVcyDVIULo/f98Phu7fi5VlEJwVXLgvLQKVZ64voi1UnfMHOugaJLKkFht+Y50Q
88rmX4Ku5QntpgJQRSsr9Lj3F8Jvw5mnyiezvxz/hEYJ2oqV8tdIM8BqeP7ZvIxD
CdpE9WOYWxdE8gnD+7ueofC2MKy8i5t0WEIjcIZCjYHTkQwpu32sB7zBcoAWcRNL
YZMwZqgxA2L+WxVcMY9/7j2vQpEXFiuM/TujqWGLjI9fKhmpDXjRRMeM793uGktw
QN4FfgVPqIf2qRqZtdduJo4m1mD0KxmW3soamc46elthJc5NxI8Pq7v2T2jLsNwT
NnijJZzM1ojpm91SUgYJNR6OEo8sKdreZhfbmXgEaqinm6ttkkahk8CvYcybstj6
K07lfacnp6z8fUd71RcLYHQN+eNQ8qEldQ2RrI9PrWTfZ7BxdgpOWcsNLfs6Qev5
s4RwuLdoRkz6t2weWdCdumSTBMPjRNGCVxlRAFW6jxTiQzTTeDEM0ZyrSgkpxlaS
yzH19O8Ni0Zq3uKZDcixI1d7k7Du9MULlmMl82TdCNh/zaIkWapnGLUKT4Sc3h6X
623yB890Z8e7Br9bwqYyLoIL76nwsoZq5npCiLR8dGe7/SRl3kt1qJgaxyNbo/9L
gdTZzsb9K9xWxGvLqr0GZ6mnjOLLP0HCJVDLLkG2gYROPjlxm4SDrCLLSBJHUcZ0
5kgxZSJeEoqADplX0oJMhXZV1+J8k8MLyF6Hd+uBT/LMv42+M2lYmu8gYs86Mosk
q5QZDLJiXjH9mzpuLbJ42hBFoT5cEtMBWLvr0I4CMA3EzXDOhIgxK+c6ObbdBGz0
30NL18LSEHm3lLmGvoGmHiI706vxzcnZ4iEhclN15aGJrnyEgx+8I57bED0q+T4V
W9VVJOjVv8+SvdyS8LU/qaqcCTg8e6kGhfWYat9A3Rq4nd9gQv9OKrLYxRUH754U
a06a7GTVVcagbr8cgnxjQFdmC8zLH/0V28R+w93+9oPuhFuNWMsuRgffGPjBOToe
7rQ16Qsp00LkORHC4sZmcH+gixNhS9zlfw9QnMYCArgAsKmUnNE8l1gNLuWcYxmj
fdmvHn5a4FU/vVPEOBKzLUGZ4TDxtmYwYCZEEcqdNYkyt13Z5jjfur0TjEJ1mFI/
JJdW2YrAygxCIu+RHeNe0HNvZQ78CC9RQSgEWWNN1DKFL2J4RQAJ+Qi+fqEx5zkB
pxczszIaVhKMcfDJNb492gWD/oV4fu0SrYbHH1aqETChGkgxCF3jY2zgDp2s8fPP
NUhQ7pbfU0wMwX6NxLajiJo1p18ZWsqsbqIIbInyqAnmWS/4psjnFGCa/WQTh8Rn
NYzpr/R1jRtt18p7c0jQCWMGHSDehn5Uju4Gmij+dbc0jmJqPYp6XoujQi5ZpOPB
zvH5hZRvXGnLL9pIvlPa020QYtgwH/IpdaRMsLB2apFSdt9PJGNX8mHjTp/PjuXb
haRRkY9G8yO5cTlrOVfFvEQvKPT8ho4p8bJ6XqrLnAzUUBKnEp05MRsDrWBQVWmA
zDgjHXzUSgUVvWyXdZTQ1hrBX8wT0nB/eZzpDLHSEqq5K2KvK28joajTmB3IJPsD
dRG8Vr8mZfSb0DSVzMkLU59LjX5G6xBWTk5id7GhSr+Fyxfnp83dcGd26naCEC8K
LCIAYzhAQnImAoHSbrfLPK/kl6advKY6MH2sS+6RgO5w8LWyaZLS6A0Bs4TkkAnH
5aAQZ9RHFHGdK+j+4h6vQapsaxl3nW8Rv0rT2Rr+X5vodjiJVSoLI1MAbLpL8Gp4
gefH/Q4tg5913mWSs8u8CtSrhgaDlNw8BE5QtZ5PBjmA6CfgIOGsptsYthC/zPFJ
AqhTpfUbk3YaWUZa0gtTcRGFfzzbBOH230XaI7EPsHwk+CJ16Xr4Goya5rKzeRow
EUjeY6QE8dKT2rusX6+4dSGLFVNZDDHbFqoycqqMQlu9H71nmmLxPIUtUqYLTQIO
q2NlEOPc7nqRxyaoH+fqfwqitPrMJnlUkDShxqO3GnFZpxRVsOynh4z5JMF+7e2K
uxRnMMr7hnBcj42pl4CVPawt+1JQn5X0DaHR8iKg/VWvy+ZBuFBzj+vIW6MGsMpU
RxfC/g32Tbe2Dy3PJgkLK9XIkpn8ysjTYovs+OEQ89uLXPWdfa3bJPnkUTG5bnW6
84rCODxjT1zSYY7V+YQ5sIJjemSmmmH7ad/YOkFjPx7sHhngB3jHGeEa7af1JtXE
9P+g8DEJ4M5/ISPB2EY2ysDZeU1zyhz45JTPyW5UGgKnkNK0jNoSQX26aAI9AM7T
tJhUh7ruCgLfyWE1QAnVFvSR8Q0Xwo57jvsxXepH9hdR8Y0tCT0GO8+jmR9jEg4r
X99sFIoOVerEFS9jbuaEne+U30PUDsH9kP2LbC4f0rcOFY0YGfOSChKHT8nB7Ols
D7i9+cCTLokbWfYuN9vlEGkwKVax93KUyw1CV4TV3ZZkBbuIDYiL02CLuleJ65Xm
F63rCcs2zj5ldatv7PCelIIsaBbEOhqz7WFygx/jcEJlSU38nbXgZUNiBcwBvz2g
cYZRatfCg6vbi9XUTuSKXIdIC+2kg0lQ4sEZ+i7Ctj6Xmcy1Y25L4SnvZRTsV1Sk
o7SEgXmNSf+3uMkHvAnuC3j2yBnlkDGkAaeTy9/OIIQ2S+Pp7MNkH9vLga7KpdxV
PkBhFnQdIxwvJi2r1cLvdgq4mFGpgfhRmeTcjTEdcAUXezt1ex98DK5QlA4vimQq
gjPGv5ErLpTqfnNXhAZxfuO2AMXvalA1fsyLnrzU8q6PI+BYymObc1Xiu6qLmqHL
TcWWxRLrEkVRhgEYk8qHC+kKDLeNN1+v0VaOAU0TiaS+oHsQiVYVA7hBe1HCZOAO
9BBmWLS/XH+ZXzZCAw05iV7sVKiv5fTfSje7yhWurzzx8fzRfaAZW/vMiKXggREj
c+rKLTuRkxFPl56SI7px01UlYbmKpnsvPOu+NT7z+Und1SS47QDf01c0+MvDpUxm
eFS7YngTJJArlnfYbBZ20tRDnp+c+rLCZr+Ueqs+oz+UP4Xwn2xinXMpa2lMU8je
sDuooKCPl9fyStLLYEoaqj/nGHH6/ui6bcYtnjrrtZIRYU/oBu5LepZBuyR0mlmB
s5vTya6bsynh4GXCU0mIPwOx4j0DD1jMrJncqkoaqMmKTad3ViQIurz/p2Cqw0av
YA/qd8EvbGyufSEDs3n+gNhVZyBH8SAtvnULWdGaLbEm/6zie+Q8vchwT3Bfw7I8
NNkyKOVv43BupAM/ijMMZ0RO/xnZada7/LLFJFKaT0o0T1lQ/f10ApjAN3/kYMZ3
QYHsdNZbBMdmKzvZbD9EtUDhzOGfogBUYltQJTwSonk6gio4zCASxeegMGzMQ/x+
q3t2X4k2pFN/ryFFJ2S1tsqUursQfbgV/6RD0PgoIYwSUYX0P1uLxUMJsHd0WF2N
mkutkZ8IfirX1srLnRfNMptYKha7EO6D6/TvQrhh6a8g3iVmDF2DO7n9UFol3wSx
z/vwgkDO2Q7USkzEpQs2jmc3+ydcw8DEeOCU2jMHeVlM+YOphxqMVY7Bw0bFhz1o
XXa1K5BSn8tbPNHsvA/x9R7HFhJ4vw72TO2bzX5hepv5cQzm2VdfRzwJO5zu2ysN
hDfGvWuFF7MOmEOVtCFfEKdFRqg94hWb7Qr7TLAO4fBN0ucLqpuInjPbTTSlgsl2
rGpzOEGsnRmDxOhdISw/XodGJk4YjIRk4HPSODZcCmj6gtGqE9GQ/FAfQH+Q8ic4
uu55n4bUdhXVZ1bVoZ0KDXYTR/xSYcp0/SxH72NWp6/p+BNi92LeEqB5ZmbdZnYb
mxth+b+QRdq8dSXzRzjhuaUV7qxV7GlJfe7oZacLTGjLHoP8Ksph9A3Lw/QIS8HD
J07gM1fAoxx82+qEzDSD//6imEB1pruRwHCdB2SEdGN67twXekHFtGE63IwAjTpf
zqHD91TALbCEy3/BzjZJ6FUAv3qzreg8qJVHmBw0YfQmN7EZzDHlymdu+JKsTyHI
WiTEWuUT2we5UUbxxF5mL0QlF9HfzjdGX7bvqHWuv6PJXaGwreC3xAt7g9C7enyM
gGaynyMQ1w6bW23OZ+7n8aHxnSpjYxPPMAAWI9xaXj1JJofpncxq/6VKzKP8mrX0
3DrpobXBvVFS2LiF0LOgxhe99DvA4RbPLGu5Lq1z4DXLStlQPqi24wGMRD7MZnQc
1WLnE3V2UA5FErynJdHc3JPko42kqAZtgy3+uL1NaQlOFT/fYT1hqcsvPUNGuAD7
yKULr+ANbedkU26HXRNun69/x/2aYhYSz8UWCKKSL1HNksR44Li/YnSzdr24/6e/
BpP6CDK04tlNBkZ0yWn3u3Pl7WHH2e+RZrzxDdjHcCWIZWEeZeNSYO8zpbl4TIpy
Cqq+dVMv0O4uLDuv1adjGal4ujiAztDz8t0nMEGM4ks5N1Rv+HTE1QY8dKMpapBH
P1l0oyf0CHtfiBRsLVRn4nIi7NeETXes+P4IX6eTJADfQHiBTKUnxym+u95Y9pYg
GEw7RVU1/ccTbuDxYNfz+4qw80z1egRbEiWXZjuD/NU7Ypx2yiGhku33XmT9Y+4H
bDC3LrEVMsN+zjkXE+eqh6vmgGOVZ1lkPqKvf9WrJrlbTNOaKcBe0BgroUZYGIB1
oIaE0LK0EOu3BtlYcjQxPX+ovPnwTsxXkAsgpMNCircGcAI20PY9GrOywaOfoNHo
l+npIEEEjhwpCkQ0igjed0Sj9KY2nf3N0u8Mh86RU4PDDD41wp/AWUqnS8hBaH/t
xrIXdYTGLv8UM1c9VoMfhR6DaiWbrtIckjn89eO0W7vfOhL68punpdziOsKyhA/M
B8XRZPlHUjCdpQg2U5glnv/2DdPlr2wk+wtmTppz/WpHVbOjSQUM6vdqwzRxWUrx
SJEVq2NPFXGfSzjfjSM8ysn08VrhkmUbdP5mswM2QFtYqehmOMINHifnfzRGiWh7
G90ijcWY6muC3Bw4Ov4VTpa+d5DwmU7pK0hRF3q2oc6Tnf2FVVdWtjgPulggV982
PUVbEiX1RMcGN7AIj7UDDq7sNOH5aniHxXxk1g/M4JWJOn+I7kO4UKnLffipAzQg
dY0MzbxudbEglfAdzvJqJKzc2Tt0Q12owdp26Zk6o8Don2XRqBicO6C7A1RQMNJQ
JB/azI9E9zDUpfeUhjpyuLfgQu5cLJv5jAoEzUMXC2DS7elmaZF+ZL+HJiiZNhsz
bpwYvp2sYLR6WJR02NEdOUw2xoT+PYrm9dC1VVm03zOMhaEQ9SmEdx3uo6S4kj/9
g/WYV4KjG06qVf6VLXWW8iPiYJsIaYNLDiuK95RyFYT71kUTLv4EdbWTDfqDM6Xy
I1w+9lH1np8gpOA1QhhyVyVl2RgqBm1yolKm98+tTPJin4WyBsGQ27vJ09grWcU8
kgVDo+rHM8NJ+qlSbjnrkkUs+/HXActapuH3xPM6CjHbriusIpjOj9iK4kRKF2io
oOgSKgI9Ggi4N+HgezZGsk3awRkR5i8I9qpvH4VDQcny5HvBcMkasmGIkLknPNRX
K34YPdFyNYY6MY83TA1kYVQNTGhVYE8BPcXIjKrnS3FR5uik4b8fLLTQJ90GsTAn
vOvbebr4QY7kTv5tpPC2UeWySKpM+4IWxgL5XtQTuvU4yy/GsSAYN/je3BQpAWGQ
0WymRfcx/dsyC+Cs9kyFSmn7IwiTRKRP1bOpEq89AYKp8/nkd6o7OXUa41YEkAE7
9LXbj9861cs+kENF6Ob/8c05gMmrAPWU9/bTh3cTa+SOdThliJv3ZyzszmL/CYOL
wBxSxdQ2Lts6R3qRJUjBnZRR0i61wYM2KQJ8kyiuulYSThacp4X9xevuAg/ITpY7
MpjQCWNW69TwWN1rC1qO4dGg4+3docgXuW83/7nMj+IDRzdVVnjqQZdetElht1j6
/LtpH7/f4R2wvkD8SAdt+nPxPyjnrR+tHzdCfx4j0JZSz03SV0/dFZvEiSuhxPp5
+6IVgyL8pRqrjVs6KesatVwNEF2A5rNay604HECiTVgC/9isCB4Je9KoG+JH/X+Q
BkVzH1Bj6/AW+ZQbPEkxmpua3lZTePH8ADUczjw2oaaVGTlKokdFHxxM4o9TV2oq
uP3KrVaxtjMflgskt0XjKv170h/rJmebZFfr1MYPh1Oxp08qCsND1vadtY2ijy/+
qfGazKSpXOCHNdQf1vRw9qxJDBLUKZh0tMzTKXxU7YN0Xrt0tB4afgzcVZCTT6hM
JZXZkaCV45LAWFrB7PNSEpJHhaR0VaGVcxM36tZ9+cPZXUF2V45T57jkKFYFCEnE
M5d3RegHZjWZSYnPQYzUtOTiMnSP26smVlBaCewatUM73a1kQdMuvT95OhGT5IVU
45OhJ0UtCIGBGgVkWylMKtGOvlefLjbI90qmYZUbK6mHvUcJ8e6Mj0rasQIUXnfA
M7VsAaZOxSwivqnZs+oz7uasCCjhpUsuqBpDspffMMGTM9sCignaOSfaOp9YutCu
dcbfIKPshh/IHhtIrT2hfTs2L3X1/mSMn5V2YsR6eDMihEF1lqsV2x6GspJU236j
StzmUC1kM+Hd6YIfmqb6hkMaSSNAt0W8slfiZ+cSRvlF0uG7HgcNRrTOSuMw8zPn
YPI0D44pX7Kwz0Ch7T9kZ5kj57/SIxBw+nrBP32q+8CvWB7lNTNYnF2MicM95k5N
zcUArWy6vGAlZd+WdmOA6w9SfFZa4Ol7qfdBrlgRR8XA4RqL1FkiKKlzwOdosyHH
nVBhnl+S2f60C372MYNBIf8vmlAbF8RtoAEH7oiremP1ayD3rYvZf1Nk70IWyrks
Kr9EmX4E4rl+ph2n2WkRtVHgyPpDOHAjVRvFr77LQfR0B2z8xRRo3AdF8L1CdfLG
GPzUKfyUHxdGhDJnFN0jD0vnWx4Utwhjly6I5pB52y9Dw3DLXgIBp7XbeRKKoXzJ
GMaxpZIEpbuqqfe8kYwmEpwVH/Nwt26Loh1sddmDn+oMyxIDm+r2XMiL6AjajFya
5zae1274p+cUSPhlh0jFFxfgvSqrBLtAj3rdoDCFEcp61a1UIpFc8gCfR9zA7nMo
c2tCUW0Pl7E5+12QbkAvFEM9I/GPgpJgCpxTUtVLcDgDhYo1ZaLCJpmdrAP/zpVP
tAKeg3H8oWW8dhcOsGm3TP/d5bknEHKxUvYeSB3P7rDMQaL6ZrcIMckMb7scqNVK
q1bmFjBJU3YNZXYGRLW+FrRaIRWKt6EoG7ic9C+WNYt2a70lIQHMzXnDYaq/vsIO
vrWhAvxDQI3EYKv3h3t8+0oQSqXir5paZaXKNn1cwK6P0QCR1rDikoCZ7TlCzSu8
Qvq5coO5+aVkO1ra6fI24eeArY4/k/NcLadDnq6GX1VWDxtzLdjva/SX0K5Hw/jP
N7A6ERbMhGhEulrlC5roAbHjVWGcbeL9FKIaZ3LYn/xXcugQ4au4vHhWIDPfFZfa
Lb8nHydTk/suUw/tXxqg9DCPWjjM6anxMrW+tA9Jtw3GPk0Tlm6qmfU11PUD8xpV
Xt6xBgtQTf15uKszoxZa6tmALDg5fORN5QTzp0S8Qm+hYlt+ifKQT9bu2q9kIYTN
LakQanTI4IdBvlzGQhmZINPQYBUZgJFmL0W6S6c2JzgbNxrxOji1cf09AyEVEWpS
/RZ3RKW7seEOgfG9CGG923FSKVPsDbBZhgaDgXlXdaLX9dTrqgwWAt92bGvJM6VY
k8qh4SChVvGaQ+3GwhOpXVGRbm3v0qDXYSLAVuAKuByiH+jtGGPGX900xXhHG8n1
v1dz8BVbDzFvgG3jbj6aq5tfcEeb/zN0vY5YubJDjYo46vGHSjIfPLOYjphhD4k5
a3TVQDHspB1IfUM7CckVJ14BCairOk1JUVkxAwLsrrsKoGhzBjGEGAZbjkJSD6aP
V4YzH/aJl/S/jyBsXPyOJQP76EsOwNpA2jfxVp/Nr4bor/uTMEvXDbKF9Svzok17
QUt1G9CORN/uC7EX+MfH0ay+RG7lMH1TuIabq0v9tThn/qRB0Z2Bp7nbyM/wkl1X
VwTqaFdoY0pysYOgW/Ob10UdTcHVbPUWkFHDfjiTkhZI+8vJ1QMx6u/3DePPQk8z
51YF/yv0dzB1Jv0ufdfgdnM7wmDI2uSYhrwRUiqvRn3vjX7ZLKibg0hLXBBfDwYq
75lk7BLOrTeQRy5awqGqyjvhZS+Qt+ekkdms33FiKQfFIoFR62AKQ2buSDpiO8xp
rpyONt9oRdFRMLgO52asfNOO7BDWd/Kr8sTMxfG5KQPm5BAwohvc3NP3qR9IajSQ
jVNWoHtrKU9kKglcjgTzAjRRo/0Up2oQBnjmYA00HYTn8eGHnpORHYORJjmr6X0A
dPa3cioZIa3U3ecAtSnb8J1XyNhMuIow0p9B9ZJ3TGdgrUeymrh3ApjA0/SXX44R
ZGogtbcIr7eGw62EQQzFlZp6ArVmFcpLU5Snv6VHAgHVVu6viJ+uIKAFaGZT0JtM
0TMe+QV82x0N1ud7WsLWINVGf6p2AFVkS5IQ+fiJxN+dlMGqoDILz3aXbHCbgs+/
3GrS1ed7hLWKZ2eMXleiYZx8IuR0CMVg3ZfxF0CxpMHj2bbQ9F4/fg99P6YrA4mv
Hyq6apkOR8F+TLox/uDwfqXKzAvzcPI+92DD04WXnGnHovbOKQnb23rZP8pCE/VU
d07k7RhaSbFXLwgPFfjkiGW6rszWSxspVVpWBMkuhf7FrnAr2dPVxabivy9/JO7i
m3fGmdfeh38/4pMgqcr0ml761eJ3b6qr7Oh4Cato4C2yB9zlIK4EYZoeSEfFS1qC
1WlU+tvHliNiejnaJy3mIZFK8yOi8jtJ8w0rlvlqwqU1aSKTW8BCIt7OpUrdg3I0
NUoJg3chGJZiljFPWQ8jmuxw8hGSE8Jm32ofscpnXTwVBN6NVYN5au2NR9tdfMJH
Y1IfLsxKu1VvO+v7+ipOFR1Sp2Ez469lNBmrUg9zyTWNjdcZiNZWixQm6hyY5tcc
2NUR+5HKqdlJDZ5XyS327xiZw+b4RSdMNKcHODf9j/2oUxaw92+ESpmgh8QxyrWn
4VVMBVVhUW9Itbe/iCcAuBqkBTw06bH2r9NZuV5IRzcy1IQUfNsy+3uyGZfKdLJt
0bwpNxdeCC84lRD1UhSkQQstsDPUovNbUTcAcZqWBJiGXT5bbWkopvZ0eAeWCr8u
Ioa1HaTe52xx8e52Jp/1dm1ETbnfuhGEP2QgWjzPp8Qjk7RWpdLvKzvOiuDC8M87
wVZVNKDZ1A8ngFgcYFERHPnInjbdA4ZXIBu4FjkEp+Wvj9YBq+auVwpTyS4A4aVS
tHVYofggCyJkqQpJz9UtDgCZDi/rmYvqyaDUtMjpXIbc7LPMvZDa8hTTDU6WYuNb
eLhodX9OELD/xTubYxry+tg7E9sWkgXJUl63wb6QU9GhCJJ9RuDINnpUb7WB2zFq
oWSvV4B3N7zLzSY9oWMuYgVuTGJiVlmbdQ8/8P2Fr6dqF4BXhuXAmQLXYMpuSvvi
2yi6nkytrZ1R4sLbITpFA4PM6vv/WCgD+0DxL5vX/8NHnuOxYMyflvJ1kV2NzbhA
GfRslfAFKNAwMF3xx4zolF9s5AA8Y4O0GQvC2RmqakJLeD/ZnCjNph1VvIQEPQnf
9zVOkdEPKcgl2KHwljtrxr3ebLa0sgvvpzE2kkTcixpKfeHbSovfHnFZPmQ2IHAd
JeWKAJ4ZuA4Jr34GnrWkwoF0dGDHGYCl2hcMRpvv5ZwRT4yAjszm5Fd3Fe38hwnu
eM6zPQU+8+1TPi6vrHn6o4H1r7n5ejlSbyEQQ6vOw3pM4IkahFfW/+inkCo/RMjn
YDNw/Tj10CHW77YamAV2vnWabUeYnVyvpx3ec3vgM0waLL4uiQyR3seG0VXnRu69
D/gNjGjd8I+Q6LfuaLsRUvGHuhY4FIB0N5Lw5Qac4AtW9+vVns21gIDUCH5kdsa5
L1yoN61kZakgH5wObWB3e0cqCa9SM5SPI2MjDqCiQXvKfT6RjlixsfNtBzeMzrUD
8x8wBQwwhHFYdRZEZ8fu2i1UudFKZmD4ZNZ+W0RpacG9SPiNv+OuwnskTF2q2Zzl
J/0EFbBX/OfCOv8IgrunTugqpbA1n3c2pNAvcH6IRMHF5w8UVeNKs+f69o3sP7Fp
HrhDAfjQCG6xgrM+ddGAME9QmmiS2LFwrD2KYl04OILGvKETs6airk+L+lCdEiaz
mghu3YdRzcIjuuz4T4rLuUzzSFQTLvbVhYNXrJYEZsUpzj8p9Q5RuUG3xgwEC16R
tF6RjnqlDEI0WaNx7Jx/VJ6WALl6T7w+WFTLmLaEOaKh8W/IKqM7Q2GzyeR/RsIp
qVK+iEssGrq/cVyLQwFCvGYgbRUWopRZ0NLwMvqo+brcWtomui8nYgDp41e0/fyU
KIWDMunpX1229VPlcuhDw65cw8AfZ7Ya4QvADwjokYNO/aCvHQ8Ynf3YgCulWlha
88LlaICVIpmOUVZeVw5rTn2MSEaqwyo6xuU6eBjvnB+GUSjc/75anWnBgYLoJaiB
gxRgBRUPeLBQm8nIDmynj/Xiv3370Wd7zIN4F0S7FMT0gTOQFlmEQh5FIYJvjTuh
XkaPK1i/iNmB/y8a6t+RLC2nhWD7M9HDmCqCAOkIeS280+FuQcr1uOoI/tEUsh7W
in8wxmD7VxZ5sx/7lgy4VMj881CBePa57lo0rJSBfKLtBqFqZiJmgZ/Ohsi6m8aD
xbz0KDnj8vU1/J4eUKVJIONf6O1ZzRXDNV7pcyC81VOs5LgCOZis4MEUxk1JtJ9E
lRqdwELHfLUPI9lpTcjT8bJzJvc++/58BpuW9aeXurY3oWYkGTcm7tMEG5heJvcK
E+J2ptXmpIILGC4zu8pbfhcS+IQCUFs+I3+cj42x3iPTnTcDmJ/TrtiBtolWckox
LibJGE1wQ5iyAluiBgUR1/HujHE0xLc8QzMfDUDHSK3a2kbwRUwhOdyMtehtPCUJ
uWO2rVayvdBTZ/B4tWwwNuNPqZCVIHXlMWtcUdtBYqqLsMPrB4SniZ7l4PEDzysd
nvpoLkcIAsOt1iZqgxNM7jHpkdDffuKREGqLo2gnnC2+SEKomVkNgLOJYEpxDZ3Z
nyeiaOTZKRA7KyPn55ugYqcuRAC+SMv3A+7lJexHIFcQdXN5EA8H8hboIO0+ZnOv
+HvuLgYWPT1X4Z6MM2mJMSQVoGl8D/DxfBQyZv5wTmsjCFkG7HFdRoBw677rtrXe
dFiP3DdPrqJ1lyRcbWa8R840CtJ0pW1P4f5jm1UhM0MdUOzHUOSN8b8GIL0E1Tdk
ebI2EU9kTRj2ywt/rkTFMuRtObdt8hxD/VRCIrIsiQnkJhWRBoRBAjjVTFnqoxS1
lqxN4rC9CvD3oMsmuK0/vMRrEtskgfwliiuovV23//XH61Bqc/swF+xk5+E9UUXm
cL5MAMeHnP6onZgwZfQYlkxXI/op9/btwv/DaF/bBfa+UMHXWIYK7+QXigt2qmP6
EaEuAuMNIDglnZGZmq8FmjgOnIAG6tEMHjlEqhOsXoD1iwV3F/SdXC2vqf2V0o7J
aDdebFn1wBHaqWGHPyNhPCclkcTRMj2fYcoOqUgFHg8xf3zYPymc28zVYwV4hvcb
IMCjNK8ABlOwnZdNPPC/Ini3oGfpLembtAlYWnKA/bS9zT1UmGoMUVfOsDhPMya2
gT5/dQjHvulrzevwT8aUXC0oCv/uK5wwhZYyASJLSj0Uw3mpj1LUQ4zZEqVWjoeJ
m4vpDMhyzMK7BDwAISja2TKsiOmXhRvjHceJ9vBDIS6rYOtSaXmRIu7SmNaZchNH
CVvGlX+0ABxDAhN/N1Ds1kbrlljbYNd5fHg4L53IN5tFrAKZ3FZ0S/10ImIgoPSx
WWCM8YFlUvSyPgfFA1JfX4BcD6dK5ZfuqoYdqX89t1pj5usp61n6gYTChUUlfTdb
gG816PcBFZjpSYsqCpqzxO2nJxl8UTYBTuqaFX5mrj2389sTb2ROBNQVHds/rrFH
jO+EC/0tik+JWIDXtLDsnLNp3+qqQWmanjCxmWj7j2dIZZk1PXxFpDBgruYP2qvi
CpdymF8UI3dSAB59JPSjDO44a/4saSmvgrW5WkUO4Gtg9hqDE8cjw0HwRyi1is0L
C9bEBv+LeBocL23O+cxxSgg1Mt4SXmvd+rAs5MO5WFdYeQiCx/I1DelWpJJJOPzm
P7hiEOrGBRWXoQ2MY3bJjdLG1YCdONhAaNMzr2UXUCWoiYmkkkYoopGCBppkRrbi
QVBzuMiLSBCtp3r4ma3/XmQr7/IAn5W1pVucVoNJJ3WuAuk2ulyquylbSYToBAAY
iaDb6WnCG4m+wFZZq57pKAXTewF9TCL67nW6ApCMdPwErVKzF2q2i5zMv5tqKNfr
yJV7mMy5ggNauLl0Vv0vt1iEKkGPAPZbOBV00E3iK6bYxNGnMeVq8nuEaT2vaYcl
CmIv3aip3a+MIXJZwetA9/vwvob6RuD3YGjxnuiTrbx4j/45wGPgmWMGSNqKue0L
BubzMuJQyNrv7f9gE46/a/6otH8YJSOVv+stvsor/C+GmfBwRum337monQgcEpYB
spNImAZLdwjtteeVWXWsZzqLRyqk6v996deQwmZEQKk/yt5ZlLRPMcsf/Id/GOC3
3wsiNZmQ++Yj6zoO/O+3BZVEz/lLG8cS/owcNW47JfKNqIB/DM7dorzW4pqO0zEh
8h1ydNb///h/a6dZ2InjCdV4HUrOJWXLbuszijhyU7IpNUfURZ43wvqtYhL3rlQB
GGLJ41mfstsHhmTyCrur+Kw54Lo6Qatdv4KDUfvOY7198Okiirwp02KYEzXkXhvM
AsYpE4NOP8qUUz65oC1QL55EjwVGFB3G/ZverlajK5uySr66p/mkyZXSspnFCyhb
4tf7d5ZNN9AvE4mmPu+D9PG/FO9ZV6Ryk8yA6VKUmWSyi5z/0zuG5Ol5UDbFyHx0
FuF08eD6Z5Rj8+SbzledIoK/7ej/qQnvmlFYoEFa/5YY7zycS0yrI4XRqCYaiGFk
1sZ9cqp7Qj0z8oAVzLJvc1dMYp0426Ce7RyJ5L/wDqSxuNzvPTz98mCWSj6fZnKs
MzbandEGMhkTpJDUJFp2wSNrG7VhpZ/h8Y364OsJ7O1ab2Bp5TOBRywgKCvgymQk
GN4SHZA2+eTkHNAjwLFf0vRVRCTb1Oxw/WUstmTZzCyNHqyQ3q5siXJWiJd8oF6d
XcTT/gwBSx7EDNhuuXGqDY0NIDs3F1AecEKUdsUP33jboBzZkINsjwN4a1unc5v1
QKWciKR77egwuqMjeg0Tm2LfMPpE3sez4F+A/OTrfeLGPPH1171pRYUBYtvQlPmJ
0OjEyCAvqOoURrqxmuDiUGdR7nnteFG6C/AlzRyjL9irNPm6521oXvub6yIyxuk0
n2XjvTdauVCnTYnxrbqGwcRmhS//exS8odbAFXaC05xUNAKRHdF2OeBTyL8haSrW
Y+7GnyUywjPyxH/BkIFsGIJvpMfeEGfL0rOEKkytP1209v8bHGVXdIUBgxhUepAt
A3A0uPcVF6FkaiZTy8fAUsxejrdcumg28OaY+YiftZpKwoX0qQGvADtfzuvya+XA
J37GTn9Pr4sAXOgO6He4Nza/QelPyGHjfnyZYrtNupMBE3k4ypMRWgi1Mwmc2+V2
zc/y7a+EQb/H+9co4XgDNroSeOAV8Xa70CulKR0093NzZ4ZDYb0CYIzZY2ve6E1k
kL4sItCH7lOxQy3gYo3x2Dg2eiHQZcXFCD72DDVOyA889yz8iv7zfBtmqQCsChi4
K8poNFqM7j2tP5we2d4XufhZplSJHfgwev8yoWW/iJ6yPN27x0Vow8ErbvdrHjYy
Ea+u3ZJf6mEG3FYq1bXkUBDwgAS7htAT4OQUi74d0ENNJmsFYd/HDiJONXarVmn8
VeTOiboXjj6Mo1OiS7wS27iz/XCkTrRr+W80unfGeqxcdTX1pLmKrwsTZy0hq+FM
C/0fBZrZ55hrY76oYc3VvApb8URwrRPn6M8XuViiuPVyJb10vpVNRFxQkw3vb3J9
6795HML5gXHg7w1/TeAToeQxfABCjuq8IO1cW8RhWrRvLAPkGGlLgV55KjOlb33g
bEOYsij/42CsrsmJd0xcHh2EMKG+BOT2Mpy4p4om1W74au/ZYZkOfCbBruSVkK9b
hlucwv7z5a4+BBPAEL6ePXMuxO8qH6mL4F39iAtBJZFWs4OjF0teopHZ6bXl0fT/
0EtDIt7kDLb9G/3H8CTt9YfELpL/FTmPJQQ1wAD9lI03wBD2hEzYj6taDqTSAdk+
LOLvKb67Fs/M1Q84BU0RjDBjmBFW7m78JMp68OXFIUUkkGCVCxU6kwnuuuZH+Rqx
XA6jL4RNiwYdjMWu7nt6DEWEiDblVJA91dZfX+giY1Uup560VACJZSYxCpoiXwXR
4upoEZdGYzzJHo7QfaSnYy4dg4/REF8y1qGNAPQ6UwEQsoNfVLtL6gCL7f53oPoR
vFl/cMnzrv13lEVHNxalRxtSmQraxHETz6oW0AOjX4N5qzYWCeqB1ngpeZ8LyUUM
7B3gqdwZf2/wZzoWMgDArqDCde1EdTxbyef5opGhILh9ZFvh0etC/XzKDpcA1OSW
yZ32OS6gqDpvvAlPfiXlQ9DIBKoGAcz7PC1asA4bevsn9kJ0topgfUkY+/ViUzt4
WznS21MQarLaO9kB3Kza59p1DvJQXdcrUQSKod7XYq93f8eMyqu5HxS1WZFgofMA
PuZTwEbXzyc3MIpy90mL8FpODYY3230L2QfDlfxuXNEdZd8q8HgxZ6U6dM7QryTP
b2/EHRTkpbxp+XevNJTY8y1C9J3dSNcE3KxgTnG8Y74ipYW2tfUCAlUAve/rHdBS
gMHElQs+d9gry6jllDcdZuPCUvkuRNOUH0+c2VESLleZHXQ1uF4qVwiNXGt/z3ps
icuti0o4u+DWePf6NrC+B1wXcr4nR7gao9+T+p0eb3Un5TCdPKvIrn+h8bAkGH0X
PmRHk6s1yC5yqs0e+yr7DZXk5vWf6ZeAk5UihZ/r0ho1j+FMi2CsLJbfxW9CYh2i
C130fLqvKogc2N179C6MLbBXoWHmht1fbW/rvsbSU8KKCZGf36CSi+wST/Vk0cZz
kAKb8O0A1CEQYgSdFsZrEQ0DW0/71GbqeS0rYc7P624u7bBh1lWVQqB+C83m9Y3t
qsTZfqzqq95AY+GMHvj5/i9zQzEaqKl24PHYFFijkuN7ExQ3nIvCaWeqBs/98w99
p4VfMx+oGa765RxP9eTQd7rq7OSFzF8MQn0qxngv+Yoiyqonl/NY00g5wMbFjnur
1YyyBwvbKfiXfvFFfWKJ//C8JccdvHgkfm26FSuF5XN9VJWdaKB6QxB/dIWRWTKV
jVWFXN3BB6KQuOJ4eB/BL4EeyCEV+24v60wiAkhBXw/ds6U0GUGYa5SrWQost8Ij
gbIoEiIY+JNweHur9N1CIHH4MB8IMILfAaagSTQYmBLhBBzQkXhlkQf0bcYbAnq8
U5TCpFMDQH0/j5+/YwfVuNpzHXWQ/fJVyf1EPXmxlgbAauZPP9dUJoaZFrTaGae/
3sY3mJUcuRSUbolI1xttHmcecNJ1F/XDD5cq+Z6aPcW/noJyIxUP4W9zlBwy01pc
GQu9skCQp0s0GD5t1R1ApIBlvJnB+9Rfjyv72GNJP28I44XAU0Q03soEyKCOfCIZ
s4M6Y8syZyJUOoHBJptVRPPLUxp+YSgPoyo+Iq37inl+xKsDkwlTW77Ro3UGM4Yj
y256dCSrLgzuQ3lfVts4W1ioRBszn/gYBsG6f3ZJqtkntDhC9lL1vM0wBWK+VwhI
vmOjMqWBAQNBPERTSWdYNe8bCq9DG6A4NRVKqjUCcJ3YPne/519iNNSs+U1ryTm0
L+uz9FS9IYN4usIaiV92PZoNBK7KBgaJB06U/kV6QAUpvAkMSlHR3nA8a1bwsGs+
cR8E0PbKGK0VbIIbpOLstenEx9+4H3HUfi7ENX7ThPZCCA6IJuCC0XP3DuTLGbTw
p+cw5Ontd5Hcc6f0fxSawDW/T6sTljvKhm8eih9T0tBvCV7c6B2g35EUSNUAknPh
+iSvBWTyF+SmG+yjPnWFGZUg6Q5w2gPw+twQwjD9M6nGPsL0pRcSA+Hv1vNFD2F5
uGeHZPUybtbOkKnDmyGE79QdQHRH/dyn0Z/ZMMUnHxCur2nafoSzg9aV+TRG0WbX
JaCp/e53+ZPJKibONSVW4xI+BXBEDgkrBEyohOi2mmJp/CBvANCGGfDwVCG7DmcR
Yw4Lkx5RfDr/ILgC7od8zDt5jawFi45ZJeJhyaL3TTlKJZ98vc/zn8/0NIPEbFN7
DeibrkL134wSnYoFGKNjIVHdNNvupA/dqOaWlOzDglfesqZ27+zIs6/+36I8gH6R
rIrwE4SWF+QVieZCB7RmjwlI3wFy4eMfOoWZzA1zNB4LCDYtWw6TnboObRGdYr8g
6J6VYnBWUBtEm9HZN8tpo1Rj4N0LcUDCyQ/ZcbTIVUqfliH2vJFscXxIpesEtWBL
UXMfRppKFi2x3z6fLQZbsem4KA350k6i72E5Vx/eSA6n0RUBo3uHY/ZxeZAQJulv
hKDU9tIORzJPTI+Brlx0wxsXkdfOh+dQ26CRgaFxCwVHng7C8VN6AZTcpu3ImoAq
VhEzjAmBbVs1H3PBhDBvyKAiaEZYdslnAaYw3EDUhPq+fz0iRvWC9i7dWyyBu2Et
gBX1PkK73P9VWnSMcNqkMSqlBzGggGAGUhooH74AJchF7aHw9VQ1GBYwlM4ggVj+
EGGFBUBUiIZ5T28ad6g7nLMnu/ezn3QMPs104qWg57BCWXAdcVYfYf6MMqmhF4Ww
RETPVEFUgti/lyyjiAmWhmSJw/6H1iljtamVeHmGwk8TIW0WidpYd5PlURKf0Ta1
Y9rBFBCiwr6GgoNynY0G3SK6M/FjRFzimLocyWXQg3pAiBBMzsY0wvgQ5TmdDVwb
hRXc96UM6QQSneCtyjF7AXjRVkK6uQc/6WZeQ9H3mqrsa/abD6VeBjj7OybORBPc
qnmdOALqIiKq1d6ymEfQNo/1MgRsU3zsaegnuZ69Dv/Q9+HkacjJu8bsIytr++xe
aL/LzWVx5E3Ms2QXpnNriHEKOJUei0pBSMOlTybbaFlItJUi/zpXLmL2GJ4MaIuQ
3VkcgRB00OVkFmkJFtZf2bnLlj+ToUIBboi8TIWMgFLfzcX1lseqnfBfMa8qQItU
z1e2W8txSTXbpU6MkM/hJV7gODRk46y852XvtrFCzppE5r0QA6dEehsyRBkbAiiE
gEGWP2XvHhPgd6g0puhVOJJ/3YcKysXKHeE7kLVE+VpBbVfSIrFeM0E3gKm0TGiW
ij/EFYsVEL3Ob8V2aUgi0pEpIs/eFGnKUvJOqhaW+U/07W/ua7V6YNtueI3UoOWL
eKftCzTrVV/V6/+UjyYCaTqb6ETQMx18F4ojMegD7+5r3e1UzwyGp/YIvuFn32vg
TrE+jRVA2oWbQGXgSmAfwwCwkefTk7fWmPFjiQSKFVCKWyQomrZYqkQBWccgezE5
oGP08B+ke/0KWSzHqHOo5A5iQoydM4rbqVfbq28b/dTFI2XfcpXlOvxPe3aScMvg
EmgtzcI3BAHnec9WXmSp/tR1YmgVkSZz5+0rGgNUTyTQw//pyXCyuyi8s+SlKcGP
TS28zBxKmqH9u5vUW7gyyvhzZSI1FvDHO7NOuIujz6dW1P3NM4jYyGyur/kpW7gT
hNCzJVcJuNgbwWU4jJYGi/JWPOmKeg9ERnYlYLNgJ1+34OY0jnf0P3434ODtucZT
zoo8nT57dD2eZg9+ZTDVV+X+BW1lBo8dx8jZMAyHFSNs1ebEIXYLVjTkLgDwPK+h
E6PWkKfiPmCbEjKjGYqzqAvNHTL07OXqy7727TAtE/LP+In1rM90Sl3/6pWNv/bO
atov86QFK+dK2urjkfs3IPvDQAifTbMURTFbm85ErsD0y4uwgRHOlH259lV8U/qT
/6eXVpAAP7s0o8vFpb9mDoEldx7IJJ6RE9foIQ+XLSZdeTG2say5ltDWGHb6H5rR
1AK4IkkvSPAZZUfgZVMIkW7hV228A3tDjnGYdOMLe/dwHa4e0RHMIhdK3lAPLuEj
Onwdxc75FAxSW4mJL37yvIbYZ+J4tDoCDINfQeqx3h4p2hypZXI70e6yrGRS2B2o
+XzYZh/QoO6MuWo98lhQwHTqXFV/EqaoOcnuoK8vVYegykeXpFT/c0xOihAOKIMJ
s9t/+rbz4Sb4VkNN91/U64yxWwVkvjxnfCdszphZBCx7LNBIy0K3Ihtyzwu8EgRk
nhQ/fPuK8niaEYpz2AOKlk1n2YkDC0FpS0zj3HtU3AlZYTGwFaizDsmLVVZeclGw
QyiflYs7oE3cEyKsdaMoKwIV3wYMXL2dr8XLpfc6ATJCPBuG9Rke1uRoJ/MXJqRj
gWJEwdIBv3PmA4O90fM9X1D1XFZGre5q0DIMif3FRZpGZeUJvU2K2kdtDZfqgAkn
/XPh+8L8I9jOr92t5c7blDgPXLukQfBYsu4GOhtgGlLxoV4fHBgUmyxFq1ltM601
x1cQmrTDb8u4OcUA0nQ/rSb4lnu6GfzG0rGxUfc1cXffjuf6BhGVMiBoHC9e3tof
b/x4bkFVy8YJ3ZIR+YlEKDVr1V6581XcLoAI2/O/0bnizOISaqdSqMs3dlrF0TsJ
u1KJVrs6zra4ZrTephxCrKXcIIEo8/gdjw4KUovzDtIRFzoa0fyvewGXgU2TZ79k
2YFHh57oSmOLKmO9M9QsPbazz9t3SuHJQRG1UPmjF1UGLzxFPkY5Ua+o/sJ7YkNU
Ae2spWKu66QzesJ0Lpo6J20Gj/GIkKkeFZy28/K8cqab9y0U0tYQ3x2642q7col3
BBtOpjJnk6xu6D+/odFqPVfMhVg/SkpN9erqmPMZ2e+6/3+Q0RQmoc1oPn8zgrC+
FYEFJSvQ1hfm/zh5l3zYbtlvjEr+aCNKI29iezNa7P9pns2R457N2VkV5PWmDgjJ
dSDUD4sdAiKsxa09aBZZVsQJzq5w3yvjJT/6kuU49vUu9ruRAl8nSE72Ifb8q8gH
k3fK4thzxj9UoNcePDpeT7oDNDH5L+a86wTi2t9rULPSWlOFB6vNsQvg6SkZSaVt
EACX1M9psHPNqWTbiGcy1diNiOAZ4OUvpCt37pgnUtETu6Qzwtf8CqAnzySXeW7l
gWR4O9c3hdgeM9XJEXR/Sq6z/nAiqwxWFxRi+AgI9SCvWkdECowa47ZqeNqsfQBX
vnNdQPhkSY+NcTgthX64z4F9p21Sz4e5Ipds6LWxX87HDUGwqjFxX2UMjaAFsU8b
XXagP+hQFfboNsxsGAt8hn2luoyTbWCFlu080Kfsz7ZUCxQEuXcB07vV6KxbVNKK
sWHEAF0oPhgs9KvtNARWlI25s92jMy5t3et9FMXN966Pmaw1EKgvrz9zmVJJKdfW
XCENAljZWlpZOXQyT7BULIoa0RXnr81ICMhd404yZGVzVS0Mq+2Wei8sxSxe42H9
H8S/71bhMzwoiTlIOHcpkp6PErJjK6Aur/Lq9eMXit5WqfWida++25txjbYp1VqE
eobddvMeGdMvPUocEGqWVQ6h/qCkLhC7GzNo53/Jx4r2EmZ8BGB1XNQc5hMdBE0Z
Xvhwm/M+CrcXy9e5r3c1Gg1iO+gP0v0laeObqgcojV+6vhZeKtasvRCPOUHSq4Yk
GJZUJ3O3wSOf7N3HTGxzy0rWQ5hZTOaOf/2RjEVABEW7+uoXMCxqscNI2gHEgZVS
8ziepYllL5WYCdKSh6FHHxLo64f8zEvZBEAyuM//VEGUzU8Ge5O6o9umh6p212y5
D11tmyiWHshlS8TxIzpKU4R7XEo4czbn8NKpt8q1hX64LN03s14If1Fyn/8T2k4V
wNJMKOlUPT1WZNgkST3lKykqfYeN1JXmEGAU9CpKdsXpbIGau/xE0nANnE4ERXjP
/WAbaleLBRolr3yuCvoSfKVQQo271ME+/2CkW8ftTW/Oq0lAixolPpornG9sc91a
VearQZaITNllrSNGwxlP2YVCso9S4qVqeqYeHNdrmcFlA2QP2a/QWhkTf5aYqeVu
i7D00ggrGmXeWhXwF69m76H2rlfne07U+R3XECb7+WM6UzVlm4+InVI7oJOnVegm
PeUIvqMaSYGU2/24TXqccYMNIpFccN68Io1tY1M65hGKysIvFV8eOonRQL2tFa1A
2qmZB5PFFJXRPqqSwcz3+cCQbqDYtW5+uPHii9zi2s/IipAfEATuUnUs6+AhOjq7
GiV5zDH2P4FV7FY8zMA6JBjfzKJX/ygTZDixMPaqENcBcztBHhTxw0asKUYCbHfl
AgX3D778JiVppLvrk0e3nqBrZpFD0ba3J8Yx4WBxkR82191uGCKgFNzAbh3bcHpD
BRkp0XKmVN6yqbknnHMawLeeOhtnXjiI0tVtB4/0lVtrlZAqlDHrANyJIi05XGTP
luDrwVPnnyJ9mXCrft4mj25tzPhNKsKlPk5GncCHeudTo7S3e0moMU3XZo6IIxi4
vePPVWZB/MzXFBV7ywSHjIhmFrNMInll4kT8vzon7/NBLuhG7c+bwIKVJoUQ41sG
6gIrMdtriWQttlgFuTDRdQN+W/sDkLxWUlX6Tuah24V1YQE5VzkOE+qJE8O4JxTo
TU8102Lf8K3ST3TXZEN5a/WbeJXnNIhGit5luBCSRXFuvKOrymDpan/5uF2fkvP2
aQPiqWMyoMGP/pbN88bFFvrY8BacT6uGTvVJWYFXMsDb9jyevZZNcPIeqPqyTp0W
esV8wKt0E77CXZbDgrRgqsuN2gFHOqvwSIZhS4+bvhWhD6tkLW79EpZiEtJwzgIV
JKL+hlpm5ia79ugHS334XJfyZBwBajxngiVpKP7/raKEoATW1AiJqrB6C3+doF+5
DzVZQt3ico0W5aDZkJz+powKBlsyiKITfeaOXmTmIDZ0nVfs7mVxPq8wQfh0KUcz
jN25NBLU8kfN6zdglvnJSH7emdrEh3DCk+V5p6trKziermAxAP83A5zQzBePHuO3
gf/K6Gg9M6keWsLBwYDd/iSh8ZBX2YUHpHuDinkFLerkW4UaKwu4nivi41sawiB0
pZHmmQY6rYTQjqtNapGsaO3JOuhLWodCxz+rI/pY8XHhFOBfODqV/9R/Mt/vUYzl
zvHT61qXWh7e6Dh4sGpAprK76g5IN1emGVR5wP9O3X4ariR7Kyv2prLMMG+kymkI
5vBif4xjio2/zF7059wHu3GPpbHsIZhIU6Dw9NTA0SiVnWzecLkh6oFYbfTd/00z
1/pamypURW8lAr0eQRq5D2Ie++DMPL9MGSMeu4oNyMSv9ETzhAE90owRBr1jUXA3
ECEuCbUexz0Z5n0bUCU6KjtEIDxenOWt08bJP0DxdOogHgutbfPiSMoB1fSQz3hd
1NH+iPQqKvaTLnkWRBB3FNNoJHpfEGovCBCX4joHVDYAFbxoWWlwuo0w7OCwg8Mb
1Ae2DtDOYNZyd5v9RTmkwLz9KOXbj+Tms+Zo2450FFj47CInWZ7XJMTYHiddzpEx
CCl9S7bG4KJgtfrJn9NUOGJScJRUndK4IJpIuaxNHEUc0n7BcHN6i8HTIwM1GQE8
O7l/EStk/fxk3fnPRD3LGia4T8X83dvmVjBJg286gvervcAhXIPcJgrupW+U39Vq
3UBjndT+uQkT36rTYDzj6R5LLMkeaNrwmZZXgcNhOtFWr6OVVXmNA7+SchyoIJ0h
uk/jOccpzFbO5zJpyRTBrN6N/xBIeFNy/fJDyB2aV1rzp6VCOUe/Wc+kcudngY5o
zzOtxPsiBq6do0Ssna8JWYdSpaKeAZTM5/PRJLUPANotcxvEJGD3FffowNTuCMZi
hcbIxKrbwr4nDEgmDKgxYfBcms1bM4mcsbld6yZXTt77OFJQiAFUIzLRJ5M9Hw/K
B62Gxjj18H6ROOM5d6k0FiZgYa4fB1tBQQpwFqsCvIwGOh2Dcs1B2tlq4U97nmfK
9pm0hJZn3BM4Xx9IyZ9sFrNm9D9UKPYe6mHAa5BUImVlUqBc3YFCkBFDlLQudCn4
Q6mNEcNh39UWuXxWw6WooFFLvaHQUAcDvpNCiWA0yCWSSkArZHgb8D5Ya3O7Q1ih
dsuQH3wV3ExP3aI7jmDM3i+2u6ZN1gxVD23hYCpEeoocZsPnukzl7xpKgd1O69la
rCNLd0C0OFeeQ4dbvLnMXLQ6YSPbku6ZbVsUr2NkT8Ai5FKb1ylKj+z2swjuUZuR
UV4DhqCTInSBHOEINyiX6LOkgwxqUZ2/YBfhahw3hRK03SgvuBfCW5hPLzGBayzs
AQi75HwvwtFQgRBiCvmy1zdgnmnRl4xS3MD5l0MnkUAHJsjDmWVeKIq8MwIws9uo
KZuJfdYcxYjq70992jwQds9SrUbFtijroZLYvgA9U5749hTIHl5upsuZABA5w66M
01JpjDUXmGspZT/4lMMmHwrOlmclTgU7WEaf+UrItM5nswYyJYTTcxdivJoRt7Zu
sZ5NN+7suktACywzufHFl03M5a73sZ0dZyVKWaPtPFLHzeU6nCZTz4ykdbBIueO6
+mRXb4iOZ3sCUbH2tocYSpuDkfsg4MqFHeNZMuWjFbjhfg5g//qAgl9LHKxImXcR
itN3VvjKbY1zRKaJY9IIBvzfNh+CC9lfLbr2BMmNf35BHOpvSzkL1XtpcHwzqH2I
Xl6jvbcoJ9cojIHm8DyhCNxOYlZgAemi/ADG6OlyPzAt9jhfSmgfEqgtqko/61oh
eXG6Af4a/66ncEU62UBo1TlWSVIkIAgWpHmh+GDPt8ToVwVQ45i75ZRnUssiGv5J
dWm5/Qa4oZhtaVZ9dnT/A7ay87JhoHpY/4TmBM8+3whBGCzD0Vi4xNN46xcJV5mk
RZhs+R58xQoafNoVFkh6f19WUPx1/LUK536aBh18pjPBW2/DNPExQqQnRpw/1c3j
CfWAVZjq3tWar+h03c0Zj1sQyecm0P1uK/XxE8fi6X5170/ufPQ4z8LEZmNlKFd8
ktg6sp51HKxv2qASFZeYXeFGfD2+hsqKLp5XIBXpD0Sd4oClljWG76BKx4OYgqzT
mEXlf14jNx1NGXwbTDFMU1CVkXEPAIpuZY/ww7oHsR4JjUNM2mPAeeKgoBUjg0AV
M+Q6e0r/L47ZoDsLDTzPzhajNaQ1R0XNlrK3AfXMmIrRHsi5RANiZhTu5gZvnYjL
rWRH6sWTy5mwPoLf9sd7ZkbZj7L1vovTkjz02r0VqDLZM1+Mv4agU8LTTJvDwqAm
+iAnnvxWE3ZTY77FcWM6ygrBmJN+z42ILAfeVBVOyrGhLa5cUYLOo5O5L8AiBQnI
6gzvaBS7rv9FZm5HQvMJ8/h1nkaTm1UIfX7ahCRak2irq38rFV23RDFIEwLkuD/x
FIPBytIwOYsRXTcDit6y43XM2uHCLmtP6jz3t3dA3FDpRW+3gaLhZ+4isOUrfM3/
E62H8h4k5jO2Nrq59Rfayx9KTd8OOjAx2jasgIt8ysymmhsCg1wmqHYtydoX0y3T
Uu5j5/xG2prpzKG5IGrwYMfKNgtgC5ZiSqlQ1EkOWeg1rSYbhGzCY73HxoolREE1
3uYGYYOLRN6ktJo52BU6wB80ceEJzu495Wrlt8uoeIoJNFakkXtZusJ/OzRpCc1Q
EtQ9PPlazHqrgOg0usg3s92MOwn2EvZxTAIm0YTWvd8lWLUDc+uP0ku6cIMfM+xS
MFT5gF42QT2YNP5IQUJcZWtmw9Xb8ZVcG1rzHBjaDLLv+hqTzPFJpQwl85xs3QEt
qsQ0Grhs0b1lD+7brLTMCiaiQZ12phktt35qAA1881hy5v8HMmPbgbZ4ivnU2Fw3
GNDUN1lyU3F8qGvyGJzC1Sen7yAzxTPsF+THX6pevNPwp4B3RAPEas1yzERAGkoJ
OWSc18A4QeOHietrHdVFTfg7EykV6Qmwlcw5iZtsou1ZVDs19c8CxyvoBQssBI27
ous7VjN9zWShWqLZP3MHqw1SHYq0ShjvZsN4O5/76Ou4kSgnTjwR4RauFD/ZmIyB
sDQ/il6Kwc6PuDKOHTY4iLUHXNksHPDui5yZa7BRx0xq8sRKjUrxFYlqvn0hcG9O
WyFq9DtBXP/CgthnyoiSxBbqyqMVSXaXtQL6782NiY8lxmzpV2wt2EcfuWTHnPe1
O6YCfsQDJ0G3VoSHzY1dBJISjEgk6Ha5iz/6lTu+Dc1p4SBRyXh10yq4z8sERCal
qdu7AYueguEfgQGPyYNGnxeh/G2jggtsSS+gkpI+GpT/oQhOQaguZCdxIhZCo962
bzRW51zZPIf+s9MlDg8PNFLb4qHn+Bg3cJS2pqkqeeukMRlRwf992aQgFnhn9Dtt
+3j7wL+P4idVKBiJjb41fpdHutDmfICNJiu0K+7JSxjmrbTLTeBNTuePSC5UQGM0
AUM09ChL4rU5OQsuW6rzxt72Q5FT/GvUNmtXnSHMmzceyeiIUuljIplDlVcuFYWz
Sy7qO+HZgW2Bng021i5JjoeXix59smwVNNh88ko/KQCx8EuxcyCXw/acJYpxr+6o
9t0ah9N3CIi91H5Kky6uShRgYbHaJRWwHmYLeL519FDCHNTnDiHQewx22ZkhBBze
qmv3S3fQBrsysw5TLLWMvQW9AXYDql1Ss2UYXAHSBgq+eZhBoZ/Mdu6+MvK5r/YI
KROsYJ8ZFL8FfRTokLIy6CWPwn4Gf+lOaSDg//P1WT3uDC6A9ZqTEgZAQTW9XL2p
8eebKVjUrHtHzRoNwyZ4rQAAef1NTdIhxnaioKF5lW9O0kLbfrb+xFo5az9FFvra
4/LmW6FXNoiXW8vBLp53oC4GWQ0r3/wv/4MoNuB/YzKzkgZYqXF8HYcmcv7k/i/N
SkoWQ948c1LL4iLzXPXKk9Xpo8jcyLK5twsnePdKnGY+8QwZqMnxKNOk/X9V0FgK
gDWTJfJ60QxMrzWQSwsTWkZ8HUlcsy3WRx/2AuPbPVuZnD4R3Xv+D0mpHCXFgDS4
rKXF8d4YMkXQF9T9//wv5sM88r6h9RhENByYISwyHQMoGDNMGcJosAz0OGL0+kK9
ag4R2sIGjrIp+B/thdOcr5BkxqzhysIXPq1awCGefrcu4JzV2p+MD52C7az124/k
wISUTvW6KM3QOvhbCEUczGyxzPTzeyCWuCwLHHR7N6fejOMxn6fZoVT5fBvJUTnj
Nd29WQ6Pg15MO0k9XUeaNa1JE9p2YPlmwFokpPXWIzCkXAsWxDdo0GI+r4CsKF5k
rexBA9pxQVjVDswbVPdcR1DzRFPprlYshD5hg2QhTDCYWaiQXhLyOLCP8UpZ04TS
wROPmEILTQxiIQE6VtMwk4SJ3PO5dgKtb+b59PDLJemh9Scqd7QpHJ+JMAjS5uZx
qaexiLiaU8gjMZ4YcdoCxyAqDzmWKQhaelm5Y0ewLoRVh3o8SbtuNdCFe9l1tKXR
2zAvoHQZN+Mp5clBHyf55FZuF67rF4C5aZKezVhoKUqIe2nGOO6u3JrXeKG/tLNG
DAqBTz73Flg8mgZ+dw6yyGZREFkK5S/IUgKNVeKmHaGBVpFdILSNmIh7/MKv8Shl
QsWVxVcGYhUC5wUV4tG8cOOVCUZRPmHDCaSXTXk3oc+3mmEzXAOj2zLhBUbaBq+2
HHcHQK5Ii3pSgn16Qzfll3FfNPjUSxXtpXnL3zySzcA2qIviUU9+lbyOT+STLUtr
UnJfpPjIa2Js1o08Xcg7PdQbtbjGEPbOndllQU2lxUEEevZXGalkDzBz7TdM1Xi6
1AhCkXzOt03cUTbYDMBenLReXMYjVlqYJISlXyudUnvMKczj5orxd7xljHSyhhjB
IfnE/ea0OzjSWM8o5JeG/fO8A4KcpOSPRLjk4aSXSpI3uibAr09hGu8pN3SM5HEz
SM5ZJG+dyKTs4w9KMPTGxqMwzRlkH2hmN2ys6ZGv8DNOOj277mCt4Zg9zu7oQBWr
wBcA1mebsFcZ6YjuVVIPw8SA7DjPc/Mdz1ANeIJQzqvbX9oIa4vCUyI+6daeKE+f
d5+JPfDuQJKWtSj1FNbptAa+ukxQAlqdFsDTGY6EE/D6IUtrXSYLLM9jVbggY6zE
NkH42Z+a8VRYdrudHk6WMeDqugedzm3EEUgz8v4bisenMtfqcwwodQL73afnL+iM
2Ynw2cazDuCC9HWWgKB6Gi/nLyXasW9ELxmtRJ5PB8dx2FaoqaMJjAsW2cM3Z1mS
QuZnSDL5knqTCuaXatT291S4tTjWeNb9akTTiW2V/LXUBLDczBHZhx+Bun6OBE8w
LQLAk/obfAiv1X/94P8f4ET96Z90UMbWv//rzRDOrz5YyIH3joVQzNCDqAslrKWc
zxjTOd7E1xEVT7ZLmcaBuIi9lCLg6gvxyqPX5oWpdAbYIyqCpn1m1GpRER7wZxMG
TkF5S5IlloQoI6ih9kw4uBIA7k3QCL3TFqa7eZ6qmDUFLxavOdIBeB45FKnX4ABb
uZoBgKfPiGnA08wEyIhs+/AvkV0fqhCPvITZ5pDAzCRtHDGVanTFQWrxMWUqojxg
4Z/F25Zak1vbrB7wqQDSII8uvu91G2pNv8Av9SmQHKvJ4NCi3woIRkoPMdHrCvmi
MDdHptlR64CYmyOtUVCtm1HgloYZVT4nlwptjD9/Uv4FaXClecsGd5xghkJT7kG/
jb8JLlxVIU6cd4R/isCY6pkctFfyrzsoQp8LxEre5zPMSfAUeW5CEIdtQmy9J0NT
NV0v+h39zmceUrLMy4dHN3yxGFd6jlWbu2mskBZmbm0IYlyn5/MNP5cVWQ/mRNHI
QdscE+3EsKcmnO0X205DAnPBBhpNPDGyhIbgCGEuItERrAYqcoLYmDhqhRfThu1a
ZqDnnBuiH9vJWuGXTKZpOYleX/xr2iRh8RJ1PJjgRnoz0qjSr8mmlDrkOizL8BJv
jWiDMSM4662w4QGl0n6QYtVBNMoRh9izzoRbsIAvJhU2mDG36IYNoT5mxvUEANDO
K4PR2c/zoHhMasGQ93vJZ2hsTYRMVNnN0VdqUq9UWrQSGYL7BOysJ7c8ywAo/Q+w
WjfWgYMCNMI/aqoVaTzR6mbQ6noO7bC09hdBlslCuFXGXSgPxduw/5Qi/Z49WlGN
rKwSsPmsOAegvXGl38LfoxNBolviiBxrb4VpqnDX3XtlxMLhHcpV5bCEGBCmRwUF
lbH2kwosg7+pzMwqyugbJs8LHDK5LfQjokstKP7tIIdZzBdyoC1RmpvdtaaZnQAT
XWW5q2/5vOKA6NZMKeLNfJAHPAwDQc5LeRyLn3qZ8Vn6nXpDdELGawB8eOOlIBVx
OGx+HDFrkIakZX5KuxA2i9fq3la8U7w1hcLRdlC4i6KkuXx2BL6It974feBae1bl
xQb0Z7CQCm/bSpE4P1BQETE2WfB2M39k4LatFy4TFTuyH5PeuNDmHI1Rb0AX1tNK
gHttx5AIri1HctzY6s1j4LN6r8ONgAkzmeOKBXmauMHqXFe2u3vMoF6ovjXvflXT
9x5qj5ELwj/bm1cw52zDyPCfdNxPvD+WptpVpmRCgTnIM4IkiduivngvXd9lbzQ4
uSvz2qqmXALfDl5zAkWZ20MONknLBxEi8CNE8GtGAmz0zLLQOPgMtKobhslhkqeB
dKuRarWa3f1o8JTEKhGgQP27VSJCMWPL/9AiPaeX1p8FiGOuV/3DroQjRNG3AY+O
h+lIl4YQwcamrHO0ymGjGcy1WrbCczKScA7MkXSEcvIryuEws6YgpMhjIP8ACHnL
LE40+SzzQXAUIf6feRzVZ96e6ClgVufKAU3K/4zXuUWgjOHnGz42Y/iaVWxwKuTa
o4QL3ZXsqSEXVMJZmqZxhTapwJlm8z0h9pqFlFmSmWuDiGB5mStHal7M83ZAbQsn
1S/iKG1+F1nBwUeX+/OzH8H1r192nDeOKwPzjNphyGI9PfufdnEda/Nh+zCS96yW
qW/H7jisNhB84w/H2WAhmX4+K3qCzdgR80jhgYzJUVfH9NV7kTkA53cxPaGouGKf
R41F4wE1CwUq6HtxaGqKCIYmn/TqdMlOK7ifp/OlZmwCKxO+ZKt3lBPlc22OtYzv
JEw0kuzoLagU21QMkJ6wHNxuzL6bXKboAVV21vjv3JxeasargWVYXa3xP/reNQpf
AjfXNTUmnj6pvk13rm3ZUSCiig6LP+X90GH0syxooseWHaEStCjJPySYxcCnWvnA
Q2wrWNnafmpQK02jxycOo+9pY/7RG2S+W9hiSNeGxiN2UM+QRZWXVezl3bnIn+/8
BB+QlNjoNpMUf8Jc8twsFahhFB8r0ZaHaIMpjTrl4En18K41s9wVS9y0T7KjpyfG
YsgP1dwLwYkYmcLDyMu7Bc+K2qpsAvUbe34tHbou7GtCe1fydnnQ+oZ5GSgBqvb1
bNBtVAQ6z7Gc8WfJKCMUlhcEoeNGC46QqtPFcgX0hjDdJqT545nopj5O++z8iLG1
ZJV3LHRSM62WYbf90FC1BfLkL+FcgQig6eBpR8OqWnskrPpl/fKQcCQ+5wyczCQD
WRDP/KNRxY/ICMdgbyjkxh8KbnPikLLAbCJJ7kCS9n6KRZKFiZt3dlsLqn+NKswv
88yepX9e2TKwNv4P5xgdCEniJzWI5wKQfbl2iglDqea/9lRwCBf/bySl9zh9hjvV
+2nuBbFyawScIHPnwNpIKZPW5+3bu9XJEVaenV8BGpqwL4NInxtO5/ypM+MO9rUX
TkcRGmfOo9B+kLw6vjc/OA0sjiArK+HvnBi1xZhbN2Wg56tdDADSeLIx0tfjiMg+
iRlk93WdifH4/4+uUtKd/qLZ+lo7kmdUe3JOysZiULI2gaXuhXSQOrnjh7BZ6gxt
LND4KFfNI1KESD4Ls1g+R2k3bNgBlxXoMGwADEqooWpUSflnVD1P+gi0lrF02ajV
U7iMLFNZ4IxACaz0tla0QwJw1DLJ8lqpTeYO4/oTV9Vz08Mrl/QzHl7y6HUCDtpq
x1gbeTJ1bi+HFXFeyiquZHMMBFas/wxwVlEvX1XE1PIUTF5XHfNk/+KZntaalrTN
HlJJNc8RkYSFBGa9EvDB+n7CA81ZJx2UDSnzUUy4APHD16HAQtS03Spx/mFSdZKX
L/39tKJxLUf7znCfiEnAcRf5FA74C4dSkMa4TsI7S/qwOsVTvMjj6IArozHByQEt
u12J9qw4IvNzCOPJJaPVtb6nl6fXecP6pPPmrKxJ73QpN3YGMtY2uk7vv4663WMT
B48Na9UGVQ9chZKB+aYyyZKSYzrlnuLQZB/aE7lOAVOkS32WVHLgE5eu31ouJCr5
4CZps41nYde21WyDV8gwEu+v863aeDQBwHC3YWTAyE73T5GK3j/0UkYzEZZOTSs4
pEiTUbYDOjGcg3ACIxGjs57nB5YGan4LEC3xY/XlcuRTAIdZUWADo3L971ByRG/l
s5MhtFtKcxmY3pIXUFOC13lHMeG2ZAM3LNh3+ZOU6Bd87JJEbGp7qJ0FSBtVG+O1
kaO/95lbTfH24G+EdGyPo1h1WX4f4eXik1uFWspzlpa3ZN6M1rcjJh23915w032U
3klC7x1Mx+wwax+28CD/IrM/KyK9lYDoBG0W+valS64uBnb3W1COFKRG0YhvvD2A
zKnNvUsTH0JLqLG3wp6w6Snjc12y1sznx54LI2SzHrGJHs0CnP7YVN8UrSUDpHRq
/QbIzkjboYbNPC8mcGNoG48QKFMkaco2GMBzJvHk1ToNDNbFjCNOdnZoeKQYA3A3
ibzD6BD7Aywo91pV/kGuqwXfubKhgwmwaFTUyDcr8EuXFsmpqmcWRyrcHZU+ARMK
/2XgKNaph18jT6cZplp/WW2cM+ELflWncE6rSw2iRRrtAojzUQ+AGHH8KCjc7YnG
iL7JlRGQKHMyHhnx/AcbGLtZRTAJDXvkwqqtksLc5t9kgXz2Kab17zmqCcKDURkz
VpKl3Ts4tihk3O2uJD7xj1ci+z2ouvSlm8AzkIStbB/pQOKk2kf/UV54t9kWIGY1
BJE93w4/jSY7BUozNVjL0G7pLPAAhi0cGmP5WpCEPFz+BGC80MyKEMk1fqtJGpXa
Nd4USF3QzkIL4i15sV3ITPQBnTlzQEbBA9DUO7/XlkS8PfP5dWIPhxZbVSYIduqw
xXxxXp5kR3c0Y4mNh82dXHyV3/SZQUy7/Hdh4OAfweBVSKLRSnu9cfNke4W960B2
wOvJTblt5YYj7BGV+urmk/Srdle1EhDTUxb0W3oQJQHtvtUnnPp9bukReEjB58Ph
sbRjyvab+vht64lCkuhcnoORXO1gMGVGEVpUvztbu8rMqfyLAcq6hVsLwi8976ZY
HohRIgBfmofRAF2SzF4aOas08tXW9/FcEU9wd7OcDMSxLROWpEJtFHIu4JcWq8/Q
SkYDOw8RZo9TDK3a7xXg5IGVg08fCR0nYwPryUPbRNQcgSOt+xbCtyK6vuSlrvuY
A0DiP3hkq05Plskwx9hN+prjtvx5KwUqtafyfhqZqgiwfcrO7y8+JhvJpzTebR91
YVEpJW6u1Nz/lN8J8Cpak3tB1oHHvRUaOLlayx3nDpDt2+smewrpLacY2ro8O7vt
sTnLG4ckVG8AEvhJKmnf30m/8tXFU7RaeIQV1DvcBLjVpSS54vsQz4eGjvHy+wGe
Jl2MO9K7/pZEE+d8aHqLE+YloF01XYiG5g58lEGgSv4P9MHhLgCCnUSSrDHD+8Rc
68zka+L8Gq+BMxPTiGuZPHzaRNS/hT7v/vrhFry17PiI2TG39Bvv4pkBBzipogqR
TG3i3hkOm2Xm8Whlr5KeHb2R+I084eGtPWJ9TZxpQF44zSjE9t5/kkcb7l0sLFAw
vnJ7o4fBweqNIL4465VlDVJsyaW6avq/qJQI6K4/YppFiaSfPmC3rt/pcTUXMs96
RbOj0eHvGtTH+3DANsTtQbNNXGJ4sy6zD2tpyavle+EZ27j2vAfT3mjoKIgW6qA4
4JSNsEBJv1ePH62lIRgepukVB9Y7ZWcw8U1grWeVFn7JP1TzSQXD8L69pZfYOOa4
UxcFF7isSYHceDRP+HfeZay/j18RqXiYCGObJIMFEdDDTdfyFUlPwDs72EteWA4E
n8IesotWMS1ZSGGcQC9lcREjYdiKVvueC3cFtAvE1GzrTm9dCTy+abCRGQLgb6pQ
5mlEtpv/n6xpKGaT6WtxQHxrJYZALX6CSP3KwG46oZLR5eehreZSSaCX8Y8rI/36
N54aq7BtZ7WOkgySDoBqbIIMufWyhMHxMsSkfqFa03Ghi5gGodLNTav9VptHlE8l
pg1ad+Gr8mttICuy9JtQ2Ra80meyOHrQM2N6OMzl8ocyP5HhbXwBRkMsdg/YDxIx
K/kMel4K+5EaKLpNLUCnLPj44WkE4u+sDwT3LCqp3Lck4WcNAW1RVXZuSuDlJpX/
NVJSoNSUiTVd6RBiSzryLHjRsBGEDSBjPp24MhzZyRKk1I1L4/VXSjuIKDLKBdkF
s5z8I65p639ZRWkjvWc2KrtRsEUL1tkG7nNHVshP/TUneQIu1blA7zqGcPwW5eOg
9UaqxHITcYb2cH3VGEvYJZR+o1aL4695qLOq+RSk+pznpZNhJaXir1secA1sl1L+
UYsS0X+mTrO4MdGM/5J4ASwBSG6aVMS4UiezuGChSM3Kx6Of7/XKQy54Kq8sdDc8
BlOiz/4Y2KEUuWvHovRm8i6RNwhdThLNXioPeunXsrUi9z8M4PBQGMxSlnjAAV8I
lJCZ+IR8y4Sm+dc+H59bZIdfxs2TUTWZqEbasHz3sFqqHDMYu9Hz3bbnQ4vqOQuw
C3tj7jUCtMPi2/aEB+IIWwZt4G6bo08EhNWHhAeN/jWMAwKPosbPXkaU9fmxGwAD
I56nUlplCAmWl44THxbfgWzpRQmYiCJIsIUWNPUkWuj/x3qH9bg1Jls0oZ2EHSFT
wdwVFhoAza7eNahKlDRiRbkphPqek+eDHWJ/g+lO8IeFJuP0sF34trtbTpOhTSsj
fusqzxWSKDRBvBTVdARvazQZ4/1fcS6dT5LpRbE8yS6u6I4Ds5mLq0WerMiAp3wL
IgKjwOApibnIeQ52r26AJ3CRtH/yiadvQQk6/Tm3r0UF0NnLxHHOCSxG0R9Spnov
UpAPONfgbOeNy4tmIKdFJMokpk3AwyxXhL4/pxPKVoJLGJZyWEJUC7jZyd+lHUfL
07e7htt0ke3wyUIVW9TOrTnTGxA+TTp+IfYjH/uj51GkKku8jMzwtSeVZ3RZJKQK
EQdRWLK1xHQM0p6oei5YXnuDR+fouwmSxHbI/IZuatIZQRmFTSgr6vYHP9LNdSTa
LUS8O+effVFPYtu5554iBtJZVVb18YKuGGb63EXVPda82zx4nIWabYbdsksOvzvQ
nAxJLhkV0WpidtTmTZHb0KIY0728/nKlk1vYQzsCbtz5J/kO3rwMq34LslP4fZ6b
d0LmYyeWxVI2gisftRYPJRQdmmAtLbz2CEWUKkVxvqGDyJnts+jOuyIGVN3S1WbS
sGXE2ROp6+lfn+Rc41LBBwTl3UJX/w8sjlfX4ZUpbGsrKBdAA+WnnDWFayCgecJ1
P7DKO9xlnESuOxzy+MrEfN5w95Yv/UN9qAKCCSkh/PO1A3QUBjnlL/nRltzoSRRh
RXNjTCtnQqd68v04R0w0E43TQk9J5K8lGVJ6yq7OimjBBYDDBBansHs2mYyaIyMi
Mz/fdxypU4ldNqzYaEjkfJCr7i+yEy9aWNj24Znbm88nPgg1Ov3SDO7zbkEbuK1O
ToGAP0aPpPMQBQ7rFGSs/aTLaKrQ20KOIdpzQ+SVZCSG7lejddhqUhR/ykcfpppl
bnoE1RLuV0Kf0XNxl2QKlR7sOA4vQDLbssIS35ENk5GDXmjjuSAy92uG0QB1GoBo
q4aCUp1CgVXzSHa8lCZLBx15uV1bqkLlvIo86ESQCqvpBx27ZQPGXrcgAjsskpby
XNC86E342uOgG2qMYcpYG8ul8pFQFzBfhyp+WUmaqi3D3ueq9X0Cmn5n0mHMrj8u
XiXfpQP923aBIgNLGDIb6FLFhU0cBcSn+7bfXnQI9WiS+GhhfUr1861T+evFWX+Y
PdQttNSzHbAfS7BQ0XFMCmJUJ9l7lwb3Za5NVsmeunUnPi5AYhQ2aAaCz17jDZ4G
2WHZzEnJJ8HLDHrAL2bkSm8vB/vgouB2M6VhJF0g//VidHhOBDzndd9nzjExebs4
yv2hXtFoBJ1Jxpkgssawa/IwFXPC0c/qvuXQgEbL3e/sF3rKhMYpL2BJKzXAR3A4
1pY8f7O+qWp1GKTa03/fkFqJqfBS/jBvZ4fkULJr2UuTzb/rk/2C7IQUo15DjA5K
D9PaTprbHdnE8bWgFsmbF+1LqiSALmUmG+/Wmls3D7bR8OIA/q94kR/coNZyNL/D
mhzUeMF5QYwnI7jnxE3tV4UthxfjRpFmjY39Ww/RsTPi7a3120QHal8hbEXlWfae
J5Bs/TvHsNjQocclLrGstspq5XtyPZe1EoS+hYv8FexlDO5t9x5ejS60TP6p9fdt
p9gm9uV4FPME2+D0nFOvbFj1vwYYk7loDq+oGExq3tgcuuCv/1hFgmbTVuOrZruA
wuSIja/KHk4XR/IFD5a/TyxHVoDkoV5s9EAcdfXRqUrgz3Frk25Ihkb5NjlnFR7j
xHdaheN8TaUo8I/J/SCoJIrJMaAp6+njR+YAu/Yhh3AFIhGmL31qZtL0LCCHZOFj
CPRBoe7M1cxoeJiCktnYCr3UUy8kCpYjQkN6/loLyPrJ9/bMN8O7P016+KUYdW8L
uLbSAhwdLOqt1s7VBwd6y4rVulW10GLcxTFku6xOl/wOsRtSR1oC5IWsZmxhFaBe
yRpIg9kUzdFcY4CyoPdtjUnsBwiFBXFRdF4zgxwO1hQeGOk4cgEUXlSbx8M575Jx
l/zmskwOFXdahJv+9GqNPbnICcU8vSCpV5Ow4yAggLDF4pk/y8SgrBWVej0WXw0s
YU93DMu3GVaU/xn5f/vOL1wLYhZnWroDyhCzFmLl1qJmfC5izCVeYK+PAoWJfnaj
rTkDmCiChj76/xaOAjXTy2E6OV0GleESYM6XK3mBJK+lW7JmlSw07v+VZvJRimnI
kfVHJ6T6+rjml5GUiA3h0E/H5Tc9gn7lgcVsp2F20rnLQ5UUfpWaD7l/9RwOPol0
KNllPJwRHln8n+OvC8MfeFqL4zODiiJIiYHUILd2SFXPJf5hAwXCqu0egI4Z+r/8
rnOkvehfaNW5Bl50+hAl5xbkIYffFnoxQAHbdjTuo8H5mOH5n44ZadA4SBAMKx8E
hX2m858rkolpfwpixZBfWH6YlcGx92sph975x6nQycY7KSYqqoJc3+1snRPELCLy
0hL1LyH3Hwb8w5dLQ3iN8gd2DRQLcsGVuW2zOPJI09cJ0gPIuQIFjp3yWG/rwmFD
NxpRT9nhUChHObZGHrlZ0ooFkFmO38j/azfkQ57k3H6IOJ5iu5sE2TUTuZwJUM9c
1I3VxqBHZzDOWLjlhTWA0Gw5mpf8Qm9c3WKu+QzYDkSXKBAC1zJISSPJzYWZEE/m
BHHkgANvIKICHaVDd+8j9+jow8fdkoFQ22/M8ghLMiSQ7MTLsh8bCYifIhVI5SFC
6hnpZuyTJfVeubMbXdVy6t3Rg+ctYMRPmsKWw+npwuQZ3FVdVJhwd9Yfu5+NrBL2
QOd5C4Ww+WzGh8/kcZP6XmDSxRcZjSlKMVYCDZwLLb19ujUayPswQCTMz0lesdZl
bk8WY1DXURsmVC+aP37ATdcRoExGYuti0jftiw9RVZ68DaH/H3aa8yHMZyj5jrnr
rMXovcJk3rz9df/eipoGxjR++Rib/r+08GuuFZ3VGbzMZ/RaDis/uXiP2fpfEAQ/
L1tYCJuWWpyCwc4/N9NoyRkIhdn2Mrs5nGDA7JT5EB8wVSDVzt5gWEDjZrvDym01
hY9Wh5n59opKORJJ89RnU+k0qCAzILPImCVR4z2J+h/tTOgC9lq5WP/tfT2ZQsgx
P1ejr5Mf5LLS+xEf/y16gPx48LBcJ3NSRpnQvmf071NSFWCa9yiGHE8MzogXyDQJ
/x03MgSoTMNeTzjdrH+R54z7pB5sn5WgXVyPy6qHm5dVPLtVWwsEJeaO79YcdF3e
dnNrDjnedpJh31rvc7AN47vH7morR4kzYjivyakFqn79esEJ6smNLlxLf6ibgL/E
wK5/9tVRu0gQ1LwYX/Z3oedvm7cwqAGyGYjnxDQNSa8VgPriy+7RpOssjtIg79mf
tNY3WGu61rzfwSVrmCLMjULJdB6//nnXoj7TExY4hWvnoMC7SApcjA+Q3SxWhWBA
N9De3xxufv2GvRO9aeOcBHa6hVhoS5GLaewsNd3y8QuVALs4eUaJcD0qFL8ytHzn
ZeGipPPc686LhHLAtNA/hPZ+hScCTrG3a+ISQVevP5F1Z8BtTxKL0qUvK2VaL2gU
Bc6PvqF0pFBEXhkQjDJbY550UGh1V6XBVb6n87q1m54lgxdqZkvFbeBCEm68tT0O
j4LCUhkqPkWN4qnkxImFNOabB28RWK7J5GrSs38vwfpM5pU10W1h74ejrPbAqieG
uMQUGydj2H1AEgm2Wzb5pStSWGUz92jJTHbNLGr30ADZPpHFDpZds96Gr/VBtmnV
bSaiHmoauH17m/qwfkr9UJEACfc//NUQb7b9+WBV+kRhd0+KRmAJ5yGMbOm+DxKd
OoYIEE50I1wQMEUlV4FfwAefPBt4+QGCZODh08GVO5dRFiz5JfN6chMFKuDueATR
YmqY6I54G4arai7bD5IR3GWEx8K3/LVprXNsQF+pm0Qza5f6bWBiLQ6/KFmdXfs0
HmwG9m3kwP8wiTGqeJZP9w9KJbij8THvGDlxVR7FYZhUMvdp/6qjJr1bVQh7UyVh
Wa6i3O82mNFmo4+q1fGsjUPE8arfnhc+6l2cQNplcG0lNVRxMeobab3WmWpfRz7v
dTS6Q6qvlSbHEB4uxTRW4ghe3JRjNj09s3xHTstdiTjfWAROP1lyrNKvmfb0iAP8
RtXRCn4kFVCK12JhfcQTo0Ivm+tNyKGEFg0721+mdTnZ6FaArZsByjX8KTJkAaH6
M7LjB1JmepY1RZ9wW3CDPSd+k6NEjzvqpHLk+AgBOYeXqxAxGWArtIlY77PkppGo
b0TppNjQXjTzXiDlndnRDDqMSaJU/tM+oLGyIiGSFWLjlOQNHBa8c6d/4y+pcATs
lFV6AhUvmmbySIB08uokz8LeKxcdaWxr19ldw5TS3mqRBk1UJt9u5DQKtkbffACN
rOvtwJaZqxi2VjCX2/KNhzMWoWe6JycYXKeLOh+tEz1MDdtFHghcCjhqFu2chgjN
2/uXqDevDvW7sf9vnRPrnzcbVH1SuEJiMnpNeV7g3gXKP6CjMIkTOEvtr+qs8nlv
OYCIghlqny8vNJsBfrzVkL+G9B2oWbdEH3KyIpsfALKkrNaF9W5Y1bqhKs+4cDHw
wMOyFvfGtsvLT/IhQrPEs7mPsmn9g10MUeUXfKkBIEBIxSic8EIFI3d683b9O9ff
9iBN9PKIQBg/rFZTGn8zn2UBrGFwqrGTux4fDJe5Xn9sqjZGUq2CePNoc/WHE+N0
vQhoENZkueWx2YDttOkIhM3UIT1INMVOlPbzpQjG2I5g9MhnSxfqIHYwOMUKxcBt
tiaM5TrfAXmHTL8NIsEpFWpbeZwJWI4zjAgf9iL9qXb91M6PYCTyHdnjmUfkq+d2
x1lhVD4qqbgZLtMCgZRoLeAklA8QDVgxkyhrFDFK2EkD6KZHaRYmomETtnDTSEl2
3pWX2brCTImaRAdfhRWp5M3TdS2bcpmCJ6TIzRwEHk3ELOuPuMlBeTfzXsn/tU/O
zd2VB2ZYNxRK5SoFPzSWCnWmR8s+0YvYBwowjOAExFskTk2XQso28pXnEAhqfZNb
R/SqYcJfcfy/0/l6o73mV5rGVNpqm3SxMmiSE7fuzJsp5qMZdNP9tilJS7GVY/UA
5NKXPRoXLl5429y3lCnvtR89jCmbB46V8chQ9c5UKj1OFpnba9XVSfLxaA2yxk7w
OcQNXyeHJsPBtTcH2qLPA529/iZXMYIwNXi0r2AwKwtrQHvpa9ULbk0t3xxeU/iM
RceNqyA0Qz+hNCBYCpuEb3+r0sYIJm5LrKESJfahHeG8kDKX1K8LU/8fCl1i4y8m
sP/M4HnO2but4qAo7rYQ7PJhJbgUEZZOEInImfVYd4zcl/YDKBTPuPqIoCQQhvWQ
EY+e6R6rrUyJfMbD9QLg2sEcWyk6XnQSQ0NlfighR6s7nR98pP0s+8V0QNN5Q0oK
ptmn5EbilrdY8F73Ddl4EwX2sHF/LOclghO1H7mBns6H7/1HbSxJQwi3Ic8brLO/
JQT8oPSV5CkCCeDXKhjQIvq/xk604CR6a2TlGA6BxFpCtHRdFY0OjUu0EyTTjj6z
uOvrp2UzEdR6KPnwo+ji3L8w5TrD5XjBO0rSSTwjtVvzumViFJBSh6v+URG+5hU9
DJkc2wkx9iJhWebEqJ1/gqIFH2Bfn7hYSTua3F6d1ulUQbhTwhEC2PcCVABuXZrR
7gITkWDAeEA5i1x8Z6YEeXK6H+i60ihqHMcLlGl/bgJZ3HEBL7QdpEQfaDB/GwjB
DcQ4ivLfqEbetYvFvXst9VGp9cRvOER40pZ3yULK7kL8Jm/RY8wWAcF3Sm+BomUf
rTU2KtjjatRpTcv35GurmdHiezKUVPQQT3OxKcM0jserIJ9w+iU2Zbid2lz/Zcq3
fsCoRqINQMz8MMqWOy8f4ebwrxqP1ZAxznh7nIiP60hCybveG7Bvs3Q9Wfx7r0r1
3xa1O/PQXBq3N3Ew0Nz0+sHYjM0kFWkW6hiIHsuc6dRcpczQo5Qh5mVgEumSMJST
768FysZxRd8FjJvTfmb9SrtAH5ULpADLaqGmPx/yaKA9Uky+5aF0H4b59riKQ5hx
KuthOleRIdCthvfBPeiViKYHMsyz5hqmFXLE/hby/0N74dD7rK35tnuj/bdahXiA
HvHVtE0wGtzBFejkfT5XnwV7Z+f/Qazx7TivlSCz/ICaCSMWkjw4xC0KcJ5aRN4m
K2CjD7Qg9zKXbDwFrOyKigPWYoNjlJUs2fnwVxqNpV8HbMw8ejAPRSjmbOSrxtFL
FjllaR8FJXvdVVnXGnenofxofWTLEbNi3P7YWiYaL4TvmUAEPwIP9ggu6thoO8Kj
AnZVIUa2igqjUO6OPhEaf9lBh9GSfiZ2yWbarQ5XOYmFOxOBF/BoeSvLOHelMpVH
Y81n/CFe597Qm2iGsn1h//nO18uFXCDAI8CFAjhcoZ2CFEWsoxHli6erkAKAEHU4
zCDdTIes6XRo51/bhEae5hpESn+Uyp14n+pwfbe/OwX2THO6umFkuEr4yE+069zK
v91Am+oEDJvlo+EzLeOeaOwZMx8RwFNzCpcP0dCRH4lOkHNTOU/o7JE7weIru17+
2RN+J3GQks9mlOQyeD8L7sDReVLLiTefXMVXzXOzRDN+hCXBnxGHR33XU5KgWN3D
A5eF2gYHuJkLJe+jTXKJ8ECT1Hlat5MFEUmEEzkwV0RMCeeWH39P5MECYtCTdkxp
DxeQ+vmMOCKWhuBVGzX72gjq2lCMplRawu7z0QWmmbi+q8UQRnuPmS+vfMRJ5T+x
JRWWrQ54mBUw+NMKCp+EVdC1SBZhlTWhbGpAUTrIPKZynDaUGxh4zi3XPbHjdqs6
aoGviHOL7BKhoeRuWrFGyITZU8iPU42C2jUzD2CduuCzoLlWBrNIXMjj0c//Rydt
SJNu8TSPsiX+bYFvNeWvV15OvBCWza7pR3qmnyt4woW7pPbyR9Lwn/t8bIHQD7dn
d/fx9g+r6u2M5t3gYJ0756wwfpPiyG+R1BNKIVZTNUcrJDv6hkpb7eiI1SBpNLsK
e0xvrWlsiv8egDHVjZLUYDvtFwnTZw5Z9j3HdN9Wo3QxwNFl67YNGioRlQW0+rrt
112n3TsbhxUsCDz7U+VEt8buigksdYgVtSvrlXyKnXmXvaA66IatDySwxagW+Q78
ZfiK3ySg1JF9LInAGNHkIQqCNWIuLlrP2AGTOtLx6CRCPkRpYjv/LOmtD86yzfN1
RBocNPRJPgN6hmnSOjMHv/cpljBJ8hjrSKpvuXMLpU0kYSG24AiLU774ZkbKOeQ6
FVl2muSfiM+wLEHGETmaJF1KctrM/+Duc6oPyzWNogcVrEWLSQUfHUQmjmh6EbLx
DhcnXxe4OXF5uYzJzP+rBB6Jf1oNaGrxDS1hXWYhZlK2iQ1Px3UZyayIWZxZKZD5
Mhr4UjDzR9n22lcK1SQ0Z8VWp/UmVwu0wmp9Uis9IDT1NjeZx1/eXIf6VV56Q+b0
EA6gU+VyI0v8Sk3ouj5/AZOvj5lWbK4b4uKUNQSQcArUQCRNYs5vxvFuL6MnmLSw
O3m6JhXJRZEVtLbVfHAxRk4sc1yOoFkH8GiVNNgLQRDbPYEff55vtnUT/vbc6xsW
rGZIfX030FSprhwuB/6m+DQZyf2RzA2gXJ6iORKTxG95fs/J8X4etyme+yiNZUQm
RavvOpdQtbz76v8DE9WQBqHJYBtNJrwPU2S+jydHPQQ2NjXUl3tXJifleJwmmmFn
q5UsuqaeF5NFR+eW1zNZVmk3o2ukQekIy1/s6eYJWI0cZNCW3J0x8udedpbvoVOi
hyKtDkVzggRFymRAJ2jbnu3n3naRkPvcx12J51j5tFHOCfbHmiosteLeHR0S3zsD
1rTSW7PBA/WF3VmqQTyNTXFR4LxFDqAlo9WIvzyHRcocpvhfLE2bVrYO1AYXoiHn
tRu/iZKpfZULzZosYOzFe1W9vaLxBJbPJ1MpaVHUfw4pUhKJnygnr8ucWvYiznXM
sEp+chSkSymg4MIYdNKfVG+Pqs3Zp95eudqQjWWek9rMXng93klNnXU3/UB3grbE
1e52mJ39eKG6YUvwPxbrPPtBhIhrlKsOwafMJdG74U/9pQcF9HDuLFkjE/QLHlmy
oRH0cHTQEbesBcRvcCHxyw5jU5UBFIRA10UJVb4fPfjEHDAKobZ+EBf6mBOHNegB
H8xS8bNCNC04lHUu8+3819iBxLRZuDHBfVwYHSmc3GrVNdnZ40Y7CV7Cld9/Xffb
95UaTFC8OlCsvRx/LCMXH7Oub5wajypEgqi4f4dkj649pcRtiEioJJVvCI3xJliJ
jZ5R1hJTEPQsMgcFCTYz2RpeubZu3qhV1umpFaK8QDM+RIpb6olKb7poYiitObfE
2vL56DkO16ebp5ERMbQCEcNOkK0+npqjEY+3lrKMgKwgZeD1HB9DhQ2ZUiyXXW13
hTpuXWttx7usk8lZpCTac9O1w7ly/6bMHCp4Sf8JPc/j1iAmLT7V61qYkZrZNdYT
EGaQEIrjoiobT+pc/KHX2jWlk95Xx42OQv271IMrz6UwulM6PiqqzPZdtOj1tXF9
7eVJ3tagrgW5pysHSoQMazM7GqRiyQ0Wpvq0YRVOHcS8orSAQ/h6s1owXokJNN5z
pmz9aEjd2oEBM2IZ54H81Uwt8f/3lBQ6lx54TKirpkimTg41d255JdEt0Y8nMJgk
JLjhVIgwpk5jxsCAbQ0wzgrIgLtzLeMVpPIcnrHKzDGSfsjXZt6C7VPMjfEjZUES
XFUb4mnhIy+ZDp2fz2oG3yj0qtPMOt6dNAOp159xQc8+ZiUpcX7WpMwCxzaprnYS
ZwqX7C/zMwGSEZG0TyD1ndI/wqbyo4BEYnHDLMaVQ94Q08bHggmfbrPf5MprhBAl
CEAUAKQQqlnzIL6wspeVsg8x53ZabnVoHXR1yH9zRPmzGC6eu7UgSyoWpXQ880iT
FCiLmxsrkJX6RTfx6VtWzRKquNUnofXFn2G56qxP9e+lnZvIYj0QtV0Pz+eWT5gu
8tBXyxWkttkr2iaOtx4a0ukt5JOAwL9Ivvgk4ZMfqGkBr/Z8SmaPz1fGhlNLcxG5
TjxoTn3Ts1jufsGEgS+vr9QTtDxsg5q9C26fw/G108X9w8c6hoPFJR5url0PYwqJ
3sgfrDClcy/0v+c+v53DypMBBjPXf29JqqiMJuleezdMWSrh4gmG2pWm6CPVyjHs
55WycaWG8r7y4XZ1Tx9AKPFGYVe1yXe87577TKzEIA7Xcceq1ieLFu6h0hZvjk9U
o+ODMuXOMKY64sAezYE92I4FZWuGn5km2H1TL5BII724+AitcYL6gh+pt4WWQ0u6
5rpOJZV7EddG/q1LydcLkvaVgpMX1Ac+aMJ9ZZy70CMcV4bYXPeiy3LeA7M1jDB6
NHbydsRgmIFOWsrNfX8s3sV2qsT4r1xikp4v+XqE+NBkuT8rhLC62d2hEohbBB4H
AFOiw0Yfme/xVIEVgs6J2JpsoclabkwiF+i3Nig+Um+cZfSA5vsE5dcLvoo7sbKl
9KtBs/lLHIga1OEKwq/UWyPVa0Qg2deoUhreVq3SDbQv4RDsmDmURx+3gODyUIju
LlT5H8pTz/UxALCwb3qU2wvxexEOkwt4i8gBhbxP2azCaVa6K+0MSlmjnyZRFFHB
NAviAfyztcEA/bozcwe5QVTOHb26hxkWWn7Xn9bjUrUAZN8C62ErKcjwzCy5tGpp
pxWghlQLrJvUI8AQ/kEGhmHOVcAccaBI3NdnNFqMEarv3fdBgvK/whx8Mbxxf/yk
eWAFkBmXfpbl4vtsICopJN8eR8ivpfSV3WLIkSa3PkvVBTV+5NdWh2p0Wu6E/7XA
6u+1VEM7MCbreh56Bgb/3If7g+vRWLA235IJsnCgJo4xeQQgypTKAUpvPbXt+AGx
7thPy69+Xwis5nT8K58fvjQkMGx8tBYq4g5j3OKlQrVdXKXMWVyTrbpE58IQkB0M
1d2wkI5bZhAKWikwFLp1Kblso9wX3tjHToDK0+qGxkSuUoIiobG/Tf6r/GfSSkV1
Yxnlf1632Tbl6PTekNNTjaaf6UiXIKKKlG24TWOmqYDmZ3HDuKJy8l95nKLV9Ely
Wq+IhU5p2HF8x+H2cltQxyIZo2p+YlTUTk+vOPS6JWslUK+IEqciXeYEO5dU+HYC
6/YuPVC857f2OGIVnA54TDqgzRR3eKv0+WrgrsRR5iaweC9ERwaGSNSqxh9uocEo
vJwDH4z1aewwgjjnucdBKZT/osvGyNxI92NBuVvtpXQWMDiP78UxfYZ6WZVFREtM
RPN+ssTBsunGuokwUsvXnb5OdiPjk2N6EAJ+68qoMXJrZtMMKRj75Rk+XoeOmDJq
Da7iyeA2KF+YvuUrzCwMoF0L7Y3kEAKIaeb+nOBkTCNgFayExT29gjS2zWQ0BR2N
qwtxtqcP47DRVjVkAH+WRfUGSiNcCZSrNrAD/tuNshnzhxpd9umRtE7uDROtLaUo
kp3RPqmb4sD9tsI+sl4dmsMNPDKsj3mgFGLRa7S7s76s9Rpc1qLSgBsKM7on/hJO
DurvaHGAF2cH1LCdkZF9M8UaU11LMdBjmmTxcYSQ9LdBWuNvoWmaymYZRetAF8P/
7h975s8fhqy0b1yCe524zMmJJGQ9i6AYlxXWg/SkfYQnITHzg2lMozqG87iQJ/b4
P+gl0uahuYjg6Vqe4kLW+SkrgBk2u5dWF1fRZNWdPMi9W+pwSJsOMknyKCEckU36
hrOKPH+HvzdXWOif6cxRv8MvGzG2rq/BV2SUsS0vMch/JRHP15xp/XZG9bHd23ND
hvN4P4Nrt3qwRG2zVbUMEA2m85oyaybwYZXpoDCtjV077VX8p7kMPOFE8h6CypP/
RH+EKTuqfwY4jxm/gXkQZoBis0u/IY7w/wTvlQc7ooXXUlwvyzKkP1IskRzppG0q
oSeLiQL+g3ya4sgB5bBbmXt/+QkjvEE5izhA2Au3sPCG+G6TtCdeX8/G0wobBp4Q
+Wqoyi5Azn7kwAqQ9tjKpLTiKnT+6CO1S0XRgW9B++itLYUI2R3ItMdhsvfFdA9f
IVaI10E687UJBS2RCEbTbHDh7QyX1DP5ntHrGJywYip8c4RZYNkJEFR9XxrTghqY
JuBd4gH4tmT73nPRUsrev5Zp7rjukokvDLFFYw5++R6Ib4kpTjVaZrpskwDrm44r
MLi7IkRRQbJcHMWFbcW/mxhYOVvp8VCcop51S+xXNaChyDyJPr6jBtjJZ5AeWb8J
2RA5FwmTxpRY0QXpxXRp3dPRwlQdJmuQ8aORz744xSC+BrAY90clGBGS7SdCUmLT
qUw0DmB2IUQ7ctAAdZ8YtpX9y78/tuimxtT/roErx1zfpkEg4dNEAfNO99M2U8k9
7JoAQrhB/G3W3gq1prf3VtenivFSrAZwTq6Ox1HsE0Jpnk7FecwUmsOL26D938Gg
2Qg7r1YaLUmEvspo25gl82RHKyPjryBHK51UdF4em3FW/bh3nGnfLY/pxLp1HFWw
V15eYDnU/iGPrsaGfJJjnBF3p3pIV0mwUPMaajkn0UEO4Nj/jxBu31JyLhNbNmL+
MySXfpNSCf/0alglLAbxWQWGEzh+QHwqs+dHIgoG8vPxVxYo0q/sLhjfVjC9hOHV
sIZQb0yVK4ggwzeJjyvnbdBgJCOu3oiGGrD8WTHzOSC4kBROP48MfwS5gVby5mWd
0HwX4IDU92j7Ag7KfJOTwZO5IfnzoYzIzd4C4IfSj2MkE2a8eZImGp7qTmWF2Xlw
h6FGIhPJyp89v/BXQ3U87IlL1gEq9+1DBgPZlPNrzpBP1sXY/aR+2pNzbeVROqvI
nc0slPKXMcVH+EDqiw8aSxZyvo3MH3na0XE+ogBBrBVgLHxptlx1zTHsp+aYfV9Y
/uK/eoLpPurxuO5dSpUTJDP5ZxGRzwz96+HszTwF/+6PVBFny383+vYPckiMzDVv
80KVH40J/TwZLzIe7o1HQe2sG8L1x6v3BvpCLo7s2Rx8buNcS9nfpUMXh/OHHS7R
wjDMkUKh5lJuOoekAOjP5WLYYij330a4l/RMEfHRY0/GtonpcBTjXbJLNdzn9ACb
ggaiuDe7c0chx75jbMDODZqSYh3Zgh4CUnO8yhVf7LUMCuHI1K2HJk8/7ZFJgdwA
V6FFgtMjLri4ZEiQzcnmce670MExUmrl1wLTlkItmSW/UGMxa/GAOM24ggmQpIYx
ksI8dfBhLWm6hr4IFvYjR88MZvP8BD3MZpuhv+fTRNMd7zAM33KOtZBT25d9FV2p
6d8vbhlpp2XFOduH1PmCLalRIH0DbsD9WT2zqwNp7Gpl4cLUyv/qtWYIuP71/ZBn
wf605dwfCCthaTMY/dBT2Djskafzzo0m/MCiTCuaeI624OdzAiZfUxvud0eqWpuy
99xQGTpCDS7WAeUuxWJEvbtSzr97+YrHvUjrO+b/7ClWjsyDFuxoI+UJzSFvcHKN
7ncQq4VFHMRI04Dgowm41wVGhDaMAGjMoqL4B8bMJkhGPdBTfhXwcBwlAHAEphdn
sBbFK5CXvTps3pPAEzs6zIh2mz7zAInATgvER7Eglk+XRNZ+klB67+hwwrCBrWwO
yfBMTBjsGdjfdeeGMuUVbmlti6sTqoT1L0VQphfDcIa4swAEpu9WZ1CIWP12POn9
jkG8/aNduVPxaM7ptUpdNKoRN08DmwA5NmU3g2rwzsx5p27siw39HipTK2B2DqRi
fZa52JcDHS382zSwtEIUkW7Kd1i7at6/tTmKaQsLB8kXIwflVHcZG6r6TwoIcfd0
DMYAbhRkI9RgddyOYn4KxFhKrHoTUv3Tq1Rk9Wm2BVgTiHDK3EQ86eFCVpN0Jm1U
Mk4neWYoPVtIGdH5+7pmeo5NSezCyBxTVUsdotslHK/8b+psI2Xhn+AjjyB616Kg
a7Sm3p4y5L+xd656a7Wkz6eHxcbXvMo9DD9+jsinPAe8zuvEIkvnEWKawRl8CYbY
adyyVwWd+OEMSspMjP52yZxZvU9H1IMIbf3EzmYBAEXWqbrCH6P+bnAzXT3TGG7M
exFGdxBPcvuuimcciOwQ2uIjcN+qMosXoexZEd7zD9NWyO6A49XcJkawoX78njpG
uo9ROXWiD3ViI54JSOmWEPoC60s4S1J6iAeo9+pl07a81KYeIhXMetGpwUp8yFD8
kklvR0etlaWXde6X5Jtm515NavbGQ5wjLPJQiiN4pqj0tal7mQBOoBUc2hDeqZuZ
IdHDI4qZ4Ez2iOS0LAxwteOMwxpcore29JqfnDE3xy7mB0NV6I90PDgz2c3X+ZyW
TrkErGqUBGBnumH3v0JhEOKN+aQs91eFsCvF5Z50XudaEmFFP2pnE5hqE5PYIbM+
vFjYBfhEA7NcK1aKF6cUx1Pkx+cvdE9THpR6Ew9ZvsWzY8vk2mmw1ZmYk0HJfQak
UuyGcNs0fHgw3HKQ/aCaHTUArViILf9HwVsy2UOeKOGaASWetiv/+SZMzLrThPIU
lesGaSi8GN5rQpc8I08gKzGxabF5W8rIVrXKFYURK+boLZ5/XSpVY6isLd6idjXR
AwCh3m6XuhdWyec7JMKf6zVqTM6Nt16iqz/lmcoxawu1p89nPn85SJOxiIo15Azr
Umy70NCszEoNDfqhwEF0MXedFNxml6ETGbyEgwqzl4Ou3VTE5+HD22oCeq6BZjyU
AMAPtjjFuJBGt/vc6PfVifN7zgd1vZBogaqv/YkG+aFIBgekdqNmzxTsJvX5681L
PZfneC5Sk9nY7fGFQLa+uUsfa2CerM4RK083SxBcsyb2Nimu6ixPmGHO6ErEOn2F
qtyW/lpGLJMF3ulhOWreJrQIfuNeUN66vF5h6ky91BD3yboYB62DzZMQfZClI6Cw
h6VPUpo0w47cPZ/vkxCm7xvw/4W60KkjqsUDO5E12mwgyBjhKVjGhFq1THqhaBEt
+CAD3YEZiWS96w49AAkYVoISwAUqbTqfKL+uLIvJOPx0rTnFxQM2YqtCiZ6I8TDM
5wGSjQWQmk0hD5SNzMHDCsbFzuq55JIv8mH5Ty0jzkkOPj+MU0dWRTP7mgLWi7TT
0mLbMJMq++qCrG5D2XrJDC118bpJGcB/dSzOdPi4F2dQYn9uuYHjxnbBpSAYS83d
+nynvBDjrDVsftN7QFOXYkMjdWT8te8g/xjKD5k/KOG17L7+IUjkGeni32v5WeGS
5zcg6ckgYKHf+5i5KrVdsCwtDhv1zYkA6OZQHqhGThHGPQYOk3raQVY8snCCVYAW
AFPmHRChSKpTF1DMG7DwRkJSmNf9ovGVgYJMt67ZQl45KhlwqL5CRwcxlf8jQS0C
076pvYLOM31fnl69piSqv5cNYlp/AVKPwS4Y0ZDz6N8X6XaIUnAB7kPOQRsygnmO
t4uItdPrYDSQksz3ZqBWh3aA0V9Fz+y+KH7lc5W1G/Ij8IP66sM8Abrw+ZsbdWVI
i5l9CZsabK0p3zNZ84xWzqzFpL8Wk8/BAWq6rDqjwCynO85OW6ZXGMz/xCkfCKkV
VyPaYZdOsxxqtLiZH/hkHB5ggYSAfBE8mteTSTcozXTv39JP2FSXsJAk+aSYBO6u
qFROL+6X81h16vm5StTh9hhGlUNpOEDxBfVhxXuQp3YZ0qkVpdtYzHLJaGmsQYgL
dRH1uheh9tC5++9s1FZEryYEw4q3j+OYJ5FOHGRBGS/YiBTGEKHYTQtIg+NKOfZN
NFgx61g7ghO/31rhQ3MwAKcK8MB3brlqra5pnEs7At2L+XzfcRcLYrBqne0TQWE/
1n8Nt0OBCPuW+OQdgL2ga96rL/GnDuFJJm1B100G0JT0X1TQhhV+d3Uh5FKOO0G8
tihiPSh2S8Yrkup3vc4fY1EcuwPBbaTAsfKlGEht2bS35SVNaJjSne75s72/59LG
n5uPtD2k9KZzKQ3dHha+4ES79yxeI1Mw2pGQzsL2wvI7GHuWio0wGgvhNBj9UMKF
LXbW86ePmf/8Y3LUsVoVgSmeYpuTaRkckB4DlYzcbO81+tyb+GcFg8vBnXGuAQVu
guNblljuEXw0zZWZV93yWJVxcsLpllUCrAVFUhq+qHi9d1i94nE+0yBvSDyKwNBD
BFHrb8Z3ISrmeoWEMRJoBApa1MG90MQIYr7VWGoESpZ4Xlz5oOnLQByiUzvh9man
zF6UIGjBN/JgQa70ucXwnNljzYIBKE9nw+RTNqU3VoZzwf8f8SpP3umvfMawrdCz
udQlZ6IiQwjEILodkYuKTPbyJQ924x8RcZkzTpm6Gt7JfpXb39TLhVoeF8xAK5XB
kOGNu9T6eBdYccY9HoP4KoPJSSJUN51rDurQEkNPXZMosz6NQZiZ6vMm7pBgeUjX
biSIWgFt4a55PUE9fomZ0ooNt8Ax+Omg8r/sp+Gw98uNIWssm1hDVRD5l1QLuOsE
UIpR7Zty5AASj5TxtT6dzg+eU/xDtMCrrqMlu8bnK4H+0Dvgm1jw9w9ND/5vYqZz
gSVFqeQHCSwf/G04CNF4B9gyepbLz5Wvh4EF/U1EkvcivtqxDu9aExZ5k3zd0rmj
AxGBy9wgDn/U9EeoPbJnuVHFomS9b+8auGfCD92ISQn8br5t8bSeM1xjaY6S5AKD
GQGBikJ57/4DvTgFCmDZ4fMGo2Yn/iyA29rUHyRRHrNN5DmJn4BTFxj7GjEReyr6
B3YEe0SXAb//Fp+DaS2NJrqYLn0V1fBnP+rE/NeX6jkXOPBs+Ux3tkGTDTzLeEyC
phFfsgG7wmAPWPLRfuUWqhbCjqFW1B55z6myRxj8uUwAUAVrJZZcmQ2VJF/nGVIo
UvCIB7GTLdKs0ORqFXc4/Bt4kRVziFFyJQpjly2b1uCbCJq7neE00SCnAwLAVKiD
nQq7cbPg74t1N0SULfF96AQWQ5yeUqNtyEpHDTGUXXuHVh9Uij0X2s28G3FqpNDD
WpZr9l5sSzbGwISQQNANFoVo2JLxEXEpTt1GAsR8lcFi1LOmYTYp4TXEwZr+EUhZ
4ABvfnuh6AIVHSeS2UHeIboHtWylRluf2FuYb5j5jAX3NelChit1PnyOFgkycWr3
6SUfyPR8Hzg7cqx6BT9W3it3izf3BUK746LDAD3kNNl+vRLGtvCq8jcrbuazblXb
1Euz8ffhducM9ECUQVnEBr3Jun8dyLDhYu3SYy5FKmK8tncL3vZZY2VQMJQ0xE+T
DFDNwOMDB7RYiF1jQ6nSM8ZrTWkYby2PXRgGh428hFrTGoxjyIrQ5eCFuKhJ7xJW
xT/X99FUK4nqpDhHraae5sZcacEL6TLInTtVJJSUaWdPrRNoiTaljtA7kqwU6ZwM
epH4RoRtFyYoepOhHWQVG6tpEmAUXP/HjGqVuhl8OIKVPJTwf0vvGUHTaf0/QQCg
Aq/pKHSeCc0g56JGugCKr61fypQvRvBLmuX1ckvZPOe9soL9TlHTR0vVQVAgLG8s
ndtb+Rf4YbcoW4IiK1ORTBKjTT29jhcAaebvUYh/zSJxYVQwYMXz5vv0l5GG/bOE
iEbq5+Z7BN35I+MEO63KfBbPTphwSKjanfEnkBVF/1wVK7H0HQybnibJ3HLabLrA
ewPOdwW4R78CCYvC0OWGBvJped3g+NQ2VnCfKbpbl+y2mUsLAdFJRf6R1Erp6nZ3
kWmH9iRERZQTOEA46ehNURcm/VufOQDhMvVIDo3rEGPyRxD4+2irdrfLh86e+KTV
HXzJawl9zyiLMzFDKO17CGDYnDGFRgB5iD+WGcBx2QyM0R4hx732d20JUKlOLLkU
zkZlZoLGQgd5djJTea8LsvtHmYWLob8712D4zxFcXRZOLMHWsXVE1xxnw3qGxOdl
WnjOlI8KcSXekFX8nfLhDnAQVCkhUeeXy3SaQD7PFDXi3qPcwrYNKwd60ZaXRr5x
JN8YqHmID7rGKb4a9gwXGu3iE6IHTWZQgzJDYw4dMzmU2rsan+yovykDAWKsGMYe
G25EPQ9opPEzzDkC3okC2qZsMR866ACGOO5AgGDVmoN2LOW837fv3rT10wMUbe1A
M819kU1jxI85Djb0Yog+XTk3W42nuPxhR7rEl6hTC0sMkwtUCLv+rMaV2qNkdnNr
dsGOd6UH/+OzElyIFspIiKXkkndfFeT4GGcaB2Qf+WA7NRmVXX+qhGjFUyddKHae
n5c0qDs4YWIiTIXunUUKU12XFvropeJ3XNxG9s4GyDwQ4f4gyshyVOHXeNGAYzWg
iW3nC+qNTr1lg+xFQ7M6jdwNjvRADdykvIeZy9W0CuSJnQBq1MtLpXZ7kE/NTwTm
hbtCze2NgI7wuoav9LM7C7oqO6HJYc7DxNk1WzgrSEg/ex2WspVqgfT3oeNanMct
6C13ixXdpwklrKhBe26Ky5ABOBva3LA2b/Fu/ubMjSOWngaau2OJIVzY4fep45VF
C9uaaASfFW5CPWB+lo3zAXffy+C/GIxRWn5ndRR7O+4xEr2dryK4a1KNRPlb3inO
Dm15Kz0M002F5GRZUzZbalaP/JGCpBzfdCtufUtcY+xwefBX7wp6EBKbLmIVvkjM
ZERDngbbvrCctSxxxUL/U0UvTZLe0KsyON8pRNlEe9dZGnTQg0Z7HuQbhCczTKyH
VoXZ6VBHMvOKQ319Kpt+h5TDfK9uXoKEANkv3eIEhtiMQsMoCIPJo9zR+BUkU8k7
oWK2exnRmtUAyHfmOrUcy85ontpnGWt/xZXW9MoG4kSPAwCTtsPFZ0h/h8BLBQ6g
9/79bjntaRSfSl3CqXOdWyodbGwyEUBG8aTHrx9nGgfm9Y76VHtAckBw3CmRGlqP
SNpi5EGjgC+K6irkbjW23EFtGJlLAHXjeC/tlFEdmd2AWBLEV3JuskeCPHdN4J1A
GWDE7GMZFLbAL+ecY5c4s4BXzfYh+9lJLFqFH6XJpBk5D7qyV/jH/+zc+2tQVAu0
fVKZXuH3GZM3/1VzoXfSuxe1dny6WFeFXhUMZkemjP2Ty9s3vYE2gLC1/ALH4hVX
UklDu0bfzD6RDWvFT1NHeBivEPiWhTymuIbpM2phpQn+LEarBhczU23j76h1z+XH
lH2xvaQnlVm4hPXoo3SG3VfMPe8ogQzrxf/dkYbPnw1jPg00VPMmwnhB7pWhlSka
u1Mfw7edEIcuQDaxfnJXv4pwE3ByaeZeaBfrKaTnEOTo6VTRmRocPdfPWRBWKpxy
zBgKcBgjq1SXm8Y57nBYjt9oMX6yKUIrd03AuI31P/Qo/JzTW8Zc6yTNd1QmLbl/
EDm7GEeD+Vi//WKUevIdqQQW2ecdeZqpq/aZ8B6ZQ+GuQK9f2YxfBKCNDMbX3f3E
dKlY3SFLSlvb1qMPRf3lsmMV3PereIwNtryoElSe/Yj1DjVfxlL2v+ZrIBfmon6J
uuzZqB69p2z50qjAbQPDSxmc8+lauHHvD/AD9n+tarlM6ZW2gCvspwQwLodmPzTO
G6eieT9bU2Usl20yq9/e3HsZTiRHns4dxnjQvIVJXXTyHoxdZnyA4cYunHsoXosN
JqgdyfyvcGIeaN8BaryIhKm4Nol8Xjo4L+p5IBl/q/C/EMu3BFhyZHm9k/jEFbFI
/v0G+CABKQmilfATvHCg3/VDFa2oKOAgrgAkrJUviliaomKNevVv8j4vUMXkGOxG
ZuRhdgpoGg3UGbryaJFy9D+Vke/wQALaeWXtIcHJjf1LFKNUHGKhs0WDRRFkphyp
Q607hIQWQ7sNu4vFJxjM5dXZEuQ6L6C7WKTv7LIaHW6LTdJb6AkHPJmUQHfNqXxc
gvHoILInuVP+ThZo5zTPizq53X8eY+/0zIbTGEQqwEjEt8bj5Yi2MjMQ0xU7kznB
plyjLdrqZi/nUQR0US1v05mGQyFtP3P0aGbBEO7i27dFwN3EMqiauvlHLct/eN/Q
CxzjxEbtb3RGH5ft5SydkQJpRdMoMfsABLGrE+rpu+Sx9P/viHH6TOqKFl5h3xtx
E9R9QMm/Fp4oaCJehrpxOWmzI1eQ9hL8/vu3Zwvr1j4UOXd2//8MMFasV3y+f+I0
/zmnHzzHasHZ6KAKlkknkw1vrLuvhv2EWq+02LtxaHKnlBTBT8k+nmwgiWlOAg6s
q+N974X27waVG7h2g964LGUfy1urBM42QkEpiypspAgH8n3EdjHS8t+xPIhN+ouZ
IkkvGLPehoPWkVeUAC3EPJhYidriPeLFJ0ysHT2Dp/X392qZN6jIVwxuuBqAugeS
GPHmDqIUSMuJWdPUcxYubmpY7i9SAhSKPtYNCN6EJfyoEsKR48PXloe92xrcPGtn
1fD1dXqDDbRmIq9YwRl6XamrETl36h3gfiLS3S1xYttCb9e5u/vk57d9quudiB0h
URHTCeC4sxWUlb8mVzJMXKoJSXvJELKP/1ym+zWLqC5sidID6nUtFsaDKWQ260xD
H06JEnjFOVpjm1lRgHsZ5rgiS220ldiY6ewBcbz+HL4Ni7AFYJjrtVjfyvmCCYgp
cnDiP324XElQtA3Zfyi6ssMAf3QG8t07o0qGXypajjqh0yU1Yprpq1yqTcWz7C6m
9egPa6kCWrHhpdlbx77IVz5kFMFRig38IMXgTZPBhZxsVcNyf0DiS9K63BMPdzhV
ctJBaQ8ObLe7c/k3tKyWADqxyrv4YOECX1m/Kj/ICqKFkZ96BVro8nD4NcP3SQ4O
yUgZYojV4vixk50o027EWyHDKKF2TO05kIM8D3DupHc8MkL4XHykFQQChbRPqV33
+fRa0ne+VecFZWZoLAm27WFSKO+XW+t9RmfvBo3jmhxGkcGHh0rvw3Mss1eGlHec
I4m615VxANZOK4lYcIVShF03Ig9WC4XSeFz+JdlsckANxCYeUE+Is8c+CdHvLfLi
+C3oqzr7EVjGW1QlV4lkQe8OF0dGuzJmdLUirUEpjW9cijqGIvXNaY2X+8wMeOAu
VTsHK4sitpzNVesF69WXr7+UNbK4yvSwaWNfqUu6g+nmLifVtIbOZ7PW61k+pczC
6eLS11YxoTRcHrgAsVgodoGXeqAphlf/+PS4zoThrutgAvJvcAMZ+w1fD18tO5Xu
pgyR+RjRldJ8AzCeHm9RwDo8F7CPX93If7UExK8BGjyMFjVw1L86mn0Gf6njswy1
YC5FAquVsd9q5L6T9WevncU4EerAYudT5A+f7dEfUu/MBU51frtmzayrdr4ZiCPn
ti1YDSMEMHhiNAEDTgZjK/2xiHVtTACvm5SyU+AEivX6aeBSyz8qHBazUVrlBSuZ
TrKKDot9wpjDZTYnvp/ySYYpVwlI1KTlf1djw+HoHpeglbOFcgTe2OZ4prJBxmTG
SdXB0BxKnjnPYv0pHwbQ450s3FyMRAY57Az0wyzr8wf0Vjo8SH/8dvwW5gKWGcFw
4WypH9Z36CmLqvelhU88wgvM1LmFLCPkycJTMFmH6xDpAPDcSL2cXaIVoCW5z72z
LFrabvIXy/2WvjxzOAVl7pjfAct7DRuW3kbGm2Y8oesxvvGC8c0kLyldQDRaBadn
Gc8p73+miC2cc/bWIP702H+Hzd5y8U70qytZ2ueomz6sI5s1guwArNozqo5Fqw5o
FmtGVM8b39ZXP+Ss4t7DjybEdtrl8nzKKnc3I/OsKikuaElu4lvSBxOd/f18UUfe
47kEfPh5sj374wQADjnehccUuB2pXVp5pJJ+G32E+vErl/7EdI6kWfjoV3fEbYc1
FGbuVBm3Ut8SR2Patkcv0rpY4AM4jxDdIsb1ydkE6AfFYhFa/hynJ1wfwW0jZj/v
9KmQLXAqhDtD3qsAmncNZUAj9yHsVKgxJVk3a4n2QYNYg2ssgX1B0T6j6ff3IG4R
hKgwlwAh3Fo6vT3F9T2Pc/77mqy++EfqlP+5IvQum5Mln31eYyMWjzIftoqdMSs1
x8hiXv/nMdSEh5fgrLoY4/b7xnCFKj4EjZiWPADZ7Dt9hbFAKbhix+OTR3zT9VDU
VdwtbhQhs1VPek+X8HeYdZ5eoG4W4nHE/C+GNe7btqZ3JixbeuQ/6hwrh6bn0FzP
nVgMPfvwsz19+EvwocUcuWmz8KQ+F7TSEX/bLNr9DxItQNCSFKJ6t4+YGNwIkvWr
pcMTXtFLzF4+/puGj8l6oFkGiav1ifXLVImfH2EiLJ1TsGApZM1bXv6drliSjuuT
jDnie13oCDEkMDyLZxW/yDqC/VOAG/Pv/qoeAKXNQSQ/hELtekjdIAPqq10DMx6m
J38Id7EugQ6EhaPp03ic9r7K+q8+D8wfkf3c2t0+0+2kqRIT1qti1vd5QSPx35KL
XcOaM3yOoaECIIs4KYs5W5iPeLuDarEE85PIVLgeMrvwF3iPbOJs7IFxmwhsoSpI
d8hoi6a43Ex7VbA/n5SqhmGhjzqmo/nhJCmRCmEkeb/rtsQtNJ9XmU3iAa5gAsxa
MTMu1tURddq2OsGotfCttlNTpu0yCWHvpZPulwxsg414nGt0KdSh9xIZwox9C98k
+KNS7GfWKXMMlbv9hdtgVJDBz6WHbX5uASIaAmcNcX1OA3zymej7z2Ws6WRyMtLw
D/ycTFOnYniAwJ/lhtrp2J39QuSQfHwIdaG9HomsqSBK3FeubNFDF/XIheiIujwg
KdKk9mdODTvJ4SdnO+OVOmfrRg0kfkFipj8qF2WunW2wMk9Hlq0680Lge0up/TGm
Ml6z7V0uI5VRdFevDhAPDmZB2rSQVKVjGGIYVGEJAHxEzPtP2kz1O0EqMCu8TP3o
PR0zh3vTRa76uzDGrlRp5kL/wadOt0Hp+rSNNMfeBYByr9IyzF6JMzxZP8ZXLGPE
BpP5WRzV2OppGSjRMBNyreACHqmuijjikC831qiwhhFEYsQBeHgaPFKvupdIHbz8
3nq6w1mp2UHg+5frOFqO7WmwzzZHaez3PYiwZstluvkZYDJTGVLM1LPyTbqgKLjJ
8TrHTKj4MfujXAkUSxSpfbxjWWwMdO49lzvguMx6n/h0pmuuig/yWkokhr59RNDJ
Q0sqi7bynn2SkFrhaa1uuCN3CMl+Vr+0dO29/1jWwY2iipSWSEI0GflLaa/ivwlt
2fF2l/M1xeK5UaLzbNHPaNrmr/yUJ59bv9C/IwVgkJrUpROMHg2zyuysn6Ixet50
3NB11njTjjbjk4SNpvXgT0LFCfVimFbSDZmDs/mzB9IpfJbVeTh0wrkbQV/dHfi+
JngjwPj6IvgKB4ENnNSRm48rd/4rOnNAjtmJTCGiEXSWsZkZvVmgyXFiQBRLK6s0
D6e4lN6tuP92+yJEnZxH+5t1P3UqpgZeUprQJ0RyIispyI2722KMKZ1Q8kbnbzKX
XV+Du1EGs2YTF1Q94UllNVT33ralVWafD8xw8QPlG+AldAUkEm3rtPJsOZc3zy9Q
GPxLEd1waL2EaZHS/rI+QMqCePNEQeRC40g74sjIbgK/oaAdbz4XwjyA2AocIibt
2+RS/du6ts/zmfiDF/F0XeFylaHFVFvtSwXHCX1455zWQrInx8u1CPXHCue2kcC/
fiUafd3hI++fyBuYKhNv02Lk8RZjwiM2TOt2vtVedyjFfZy5mhjmnqDmo4WfTegR
SH7fg3yPlS2ZvVG+7Tjr9hupff795PM3xm6/oK0ZigjjtsPfprKDsBFkYE/uIVeb
0kLvlN4nAitlqI0HaRN8Mt/9N5y4Dv6slWWFMlST8BjoO9rRALINXgoEmrGxHT29
bhlD9sQMuqMCJZptwYq+coKDLyufL+ftiw3ms7bEnydzPXnLMWQZLJGz/Bpo92vF
hDq13FVCskeFpw0df3LrrgoYsir+tr2vNv54RlbZ/yTTMXyaXOqde/ZKtDdrUGpp
GYf3cGBNGKne+geWuAJmMTcMu9MBMQnoYjfJyurrbeimhvh8D9lKxJqToplCjbyL
e/bQ9egAUGgzsUr8nHpO86PbPhbBgMl8JmH+S6rVpBNYbFv9VyjT1wgtjIzqkG1N
ybhl6EgDGUaG1SBQkWIew6myy8BUWpYUVe7Hej50XJgDn6qC79I2u3gqidVSFtY9
ZTIK+424iXixSqpRnjDkuQpNbLBbpu99jHfXU9kVYgTDUAdk9YOPRPtyA2G7fxL8
bdvCnmrIQnEz5T97i2psqCVubNg69TFZS0VuEyFUezumnsisUfw2BStFI3S/OLmR
3JiabGc6MmqaGWZz5/zbz+13A8DPj6GNL6fCKxKGFY77CqJgambB2M1fEj7OYG0Q
/T0s99WdJFblfWGI7DQ5+qiCj7BOmTdrVBqMOFwahVI0YiEir+F6+A8ARRo6sCxD
7OpAnH1cks4NaarxCHeGWc/zElmAE7Syd1PaJ09PmOGToOGis5UVueR0+k04pI4i
cl/xd+ElhTWrhYP2IT0Q0xqQdZv35xAUM/4LE6v4x2p1iJudFWr5OMqFfAhh9Iir
LY1SOsUdTzISS3vm5PF8RGtez2KAJMH9wNBW2VvAhNJslOBlQeI5n/CnjqpdoAXK
9B2zibWiJTXDZBTxvy4AWdh/FVhZHYNKqNG2ji5wIElH1HkpvzdG3LqoI7YENBc0
0AoBKv0YLudi+BQkA3TIQMALDooZPB7dGJyP5+UD7chuq2I2p797ualhCeqndtqM
QTcEbZXGzB4GB0KJr+jVOz1XigYJoSc4Bcgx1+FW80Th6T4EVgoqBcOoWPsxDbZe
rqMDrVkynStyD73w+v4garGxAssKJZgHSKd8wm0Yy1AfU4lvhULpMl+lu24rTPcZ
tjEy0FMgp4lfOneGvYVzko8PUybK64tVnJILIrubkfP1+N8qolclAHbu3ED8BXng
QtdWg0ba29za9BnXLVFDDGm+6TWDeSdc2i/cbHW+iLX/0cwk/oUanBVGvt6Rmo6B
7ql9xBLCAzRoYlUp0TqSWrFcC18D2kZIjdVq2CTMkTgMx71i/OAF07DrgCyWGDGI
OKNsOyef1lL3d4DaplwI/xK294riQcJnthsz4i89v1KxU/3HFe2JkzZTgt70pBlB
zZzncRGkY1Y46ei/Bt3SLauhnF2q7LwSg9ZgGQ/nb+df8Vb+Tq8xX2RviYHmxLCk
GrPawR6Bn+R9ut2j4ayIPpjWjFf/Nwnw3eeg/s3S1vxYKhZayvpGWXQQAwqE3N5W
uendsCPxzu31YMQghCPchcP2oaQpHOWYYGkqPdRR8nTIkSQo0dUrC95y4H7wh2Xx
VKNPyljjt3X3CGy+aVN8b06FlwdNhL4iEwU/xp0Bd5tZPexUOftZnfeMVGfPTBnJ
xoo5ZUoaxIwhEBbLphzDur/+jcEh+HAHJXf1p1CnlZPqKF2aPrO6nFAALlvsfB5l
Ox+jQH6+aYAkMJniDQNt4g6Ml9t8RSvbCSPyhQ4RC0dEPIKw/w0mSv1F4VbCpdXk
14b1In0IVtwIRvCpSAEnVTqhbudcV8vhkR1/2ici7CsbwXYMmywOdFOUCack5v5D
W/G9hTzxCC7iVsMdQVki6f8ol2B2+LHKPlsHWDngAJlgB37pmvg+SqxkiMw6snda
Or5q0qu14q5ZXqH5vlDHbBCQCF7F4YpTGeeI6dO36IYevmje4ZqIeJeaPm+ocY12
5yK1ZzBYLQ7Hy9pwVuarNz6AXzuED6RUgDEX1l5YgV5lL9wYHPbfnS4mAFAcDVsq
XruOg8Y3wIIzN8nRLO9MRQ9cEsPOAASyQqRx+zWnKfZm0jDMlL+FMI7Cni6rXnvi
qaK1B6SadYf7573w+0L8goa6b5nQiNntPRL3x2i1BRkQ7eHrYKs3//6K8X/WKMtf
IRuNXhRmzGimIvPvS1DxLBaTzomE/D1+iGT9xbQbZamq655AMFj7QdT9vtDBdnm1
3KO5/BuDYp4IFO8ZkckATaooPyGreASB0yLu2vGzt3H0jUMGpFABGVPQqzuiCjis
iQTM/jXmDkN08ZYWGaqdgmeeyva0RiGS8cGhIe2X/CN6wMYK6F0iWge76xRSP92r
1bzvO+qrk+aj6BW/+i+wFTtT3QEi2qz0DcfYgt4FJPBj1DKKi4MFX6I0UnlQtma/
CPNTfFA47GLgEEb32J9Lp/AK2b3mtCRnjbXNYihhEq7vIY64/Ar6MQ8pfvLevVt1
vBMkHyn3uNC2gpbkRgjtHeIKPv2gMQinHPjPGM0XoTXHE7M3CaqXCRVaS9fxesaS
Vph/hwpL9JvL1Vqbhr/9tMuAWv2cv+RGL6TUM8g/VDoWkBUfOvzFwfBOGxJTt6KV
X6cfEYn8HAwi2C+YayBdiYchkOjs4/+ttCyIdQlAiYNN5TiVyU/lgIMjCTlappLt
s7ZM9sUuh/n+PgJUv0JRsBzS6FnoYbnvTtnBP0XRozIVnzP40LfJMNus5mgsbrrW
6weIps9dtUb7PphRDSsh3CN4UTxSNnirGxbPV8nTdan4brBu90w5wqPBOIS5IS+z
T+ZvPhxFNh+soZMcdIIeESnwJncQB2868zqYW2B8bMWxBpztD7ydMKfAwJUait+b
BE1X0CXvAurWU+C3xfmHrnycYmgpvmDExnT1jXbL1s5YL6sfSvnexcqhd6FNwrBY
se9q8L6fDrSdpFANvLaYwUHOpQuV4M5oDe9IS4KRQnP2C2XMjVcs1Yh2L5vW0gaX
4EWBrRJH7QOCliXzW3Gc2O2kydDMjC2Y2mzNseIG/NPQqaNeEgASIYPI5+aIyc8j
m+eSrSLw6DYn0/aG016DZwCK5AJJiCqkM+AqrpzuTe9V1A8F6mR0ITGEq7jBMtkl
kl7DonzgmvOZ0J7gN8R4E5gR3dL99ts4jIEmELWv2aYNC3POY4+HW2xskbGcBr4w
LiC6BgFwvjjUBZ5MYkEPi99k5gsrUFDJwds036RJH7Xm3GlqiMQv+qD5aVC6Qfv1
0baO1q+MH/obuMhwjskE0Ad3KV4PDIxcmKXfrxADdV2oyXzmY2a/9+HoBzAYKCnW
unDdrr2Cfy5kptvTaSMfQOe1csS48uF4K0C89VzdssAEdI8g7qqZ/Oee3qLqOnZj
Qq406OloH/dsTyLzLkGuBYRk7MHUrMVilXFDCVhB0Z64GdWzdRwX3iwxU8araXo1
0/xowpZ9Ocpwe6H4VS5vtVYrWGSi0btE02lEfPDB7ty6LdqfewN6ivAIySGe5tfj
1QWwwCaiMaKZTZkfREgwbDeWP2YmoCihxP/MKwG2LubbwfICl5TaHfYDbQ0QgTjM
buPvCO8l+AvQX0RHzjgP0SZR/hkbBJZxDIcMOS0c6Kn5YtTF71GD39TDQ2DwSa0m
0HbX/DpayiEGXzOhA4Xeo5THQjbR8m5PBhdlDhJVB3oXyNaNS6bxRtoBE77OjRYC
opu6BaVdGYDF0XRUwN2v/lGYxNG7l8j/prW2WPgS1RcmMccqKBXqfm/YEtTXfZJy
Cg1X+lCwgWnIGoO6zP4EBf7CLn09E7bXeOTzRifD8fnYh/3DFM//bntLEZ0qrl7g
wkO4bKo8SIntE7LnyGtZ+A+2+nyTjWFb6fcqNPR19KpTrsnWlZnEPbc16Xvd01K/
w1IFJ6d53eBKwcEWEaty9ZgTdLjmPYt8TZzRJlwrwqIXJyY4HY/2yX/RbuR8o4CP
Bs2CVlgCAXEYreM68UWRIdancZIN9DpgFTrU7MudRvInIPPpkyLwOp+fir8sSdJ9
kSWSvxOH8VJ2rp2qqXj8KiQ4KEPnXCv4uEQAkCNsrvfIlGpm1T4fDVbGJBEoFdYJ
8YMjiT5FjRNxpa3FI2wM3DJcVYLnV3G/bIBHhfe/A1nRj/2Gmehl+U4DyzuN82YD
Cwvtv3rvPWyRBPCjHF/MKy5sr+bm17vlQ5CZvnBpVENbVRGmKyTHT9khiU9ftLcY
7/JQuFrEO4Da0J7nvxQAcizHsslky/w/PuxR78YMrjvTBr8q2tIq+SIB+ezz41Dx
vc/1zOxBTOq2htNF9W72rjq4bRWJXG2nxJW2OqyMK3rUYNg0X0yAm39Qw1ayz0u2
pBIlVd45eeoVYfOdjcv2J4kOxAPc3AgZW/2l+Yq1MR+NwIlKzibRoRQtC9shaRrj
TsweP/JwWKwnocDtCkb78h86qJAAmkvGM1cdM27sxSQVI0VDLSDVQmtwPpS4cM6S
w7dxBpQhrCA0Asao/lD+l1dTyI4hP8rsNhBA4UGhiOHlROPsHXt1C6F27KIQj0cE
ThazBDbdciL7F0OClh+NGtCGrepU2U0BNz6aSmop5Cojon9vWr8Wj8pFEi5SjxtZ
KJxo9TH3RfXKkPWb1YYjbxtxzsI1ncPQ0SDJm3ydGlOQf88ZGQT1q3PbplK2nqd6
rAkB18oydpVkaQYJCy87KIItjuDsHWo8TC+OBa5bF2KCXle9Eob/+9sIp1tRKWV0
zXbv9Ukdpe1viqlom1iFnycOlyGBkXQuxbAog5+AVoHvdK01c1Li6Ckar639NGLy
HH2qMxaPqJ2g1KVeUW37uB4yV61h4SVtERoZvEen7t0lD7U3kBb3sjlAtDd+cg6A
DQDjIshlOmt24HuCPN3fT4IyC+9TjKiYhr/XZulRyLvXokpsTbM414D41W+5P9vl
HD+YG6qTf7JQVhux9BA4nnGTJGK0RPzcXEfN/7LyrkJXRK0tKaZjT6Aj+22u2BYp
a/TEPRzKfgR+jnaaFAVMGEIidTO7jUOxGufLbyIuKzOd6GPY3lK3cszAXFhXqO6+
sOnolWXmoAfYg4NyjEnr3xw+j83wBaraHQQHEnHMxmeVG0k88kzNhToKuhgWD4jU
Yew6bvkoYhJ/7paZ+m40pSqOdM7DcyhRCsSUXtOmnroH3DwbGEN1cZv5tzHqO3yl
RNfSK0s8PIYhWSS5O0Lq9Wc+lcSsMq3kLDZ3GxHW5b1aGGVWUPNkGZXmuS4TOnDY
7c0bey8FS+AAYrkkRKEhV7CldSJhTckYn1szbm6svWRk8DZ0yu6BUKwiLUJb+n51
jYwqiObqcIx2NEbwUeMFKae+RN+4z85nPDMXb92flThiASK6Z+3kx0V9kfae/2mL
UCYRumOvZTYalrzdNAXqi0p6eKUNIr0DU0+Wkwydzb8pmTb2ousjpIXGn3aD8Zux
GYp64cgAloiUGDkoSCmTbm/DvP20jKKfe2NKMEw4lDSwYMHtwQBcQ2DWVgOO5KDl
m0wKcWeoMQOubmGb6Awj0uIG+iMbWlFQgF8PgssMLPEwCi4nlyWdU0k4OwpxfkQo
PPr+ipf39wh7EFn/hOrqquJ6/auMb9mxYPlB3Nw74anu76vlpaxz2zhN/ynSJrHG
5X106+0qGgQPZ83GaVjV9yXyHhRdWNUdlxX801jIhFmuxZRYEwefEdWLoBF4mhWq
x+nsrk2Y3bogH6bnByNE+bQIVKXxM9ZfMhavIxUQFKbGo5xwXkA3NgxbWevAafFy
2dDY79Y7HKyCOk7SaF+J80FjtRz7VF3Fc7XjH1UbijReU+iV5oKZdAzAOeQ9o4wi
TMcjP3yxEHg0k3ico4U/w/C3GAoU2ZFc3La4Xog+PESCVZ/vle3viRRA+Rrqmh9J
W+4yUUQ22HZ320JyTpqOxdhO2W3bN2nEBanebAjIHtG57a4gKDmTdxn3jwJ47Dr/
JWeVGNQJrxoBB6eEoBBY2mOQkP8boIFTDxJI9tbF7Skhl2w3B6gcwZ4hULkadKQz
cL9DnH/4N9XMdAxKPCuFmPxPPZfUUXT2X+9y6fQy4l2ZzGumJKxWd2oh5tXXsXWn
esjtrRiIukj7CNMbw8UFpkeAXMdr5eut7lpqNagWJ+tj2iWJAjhYkH0wHP/3tnO7
cFrJo7W2K2yN6Cum2IEbIO4CL1Q4mqp21sMPjd7KRErJYpv6JCHHw4d4mWgllSUc
WBs5g4UMUCCVAE59+YnKXyuTS+F1kqzf2ZPuOdltdHB3pAIn/eh6JE5uf2nY+yA+
ziU1+Ofde0EiJ+KoKOs/lsYQk/i8wBQzFwL9lF8vtJsY1p6uHHGztWCOasNtSXzo
USRWq6jWVglUDQ5WttvlpqXvfSjK2W4wjH3Z8CA3pO0XtHsqq+Kn75XsMbijtWhg
HNfjfYcq2ReVmB2ZVJNaKg/kYlzKRijvqFyvdiSw3ksete8Nm4Hys8RTEfTNsYlg
Y6UQ/SmzSLkuvuDoYLM4AXwHZnoqL8CCZUCMitJET9H3+g9rMLZs9tq+YT8tlrtV
9jOQ97ixfPGYQUYqmw3wzC+PUGM2qrOINndU80stcgz/0WdyiC7AZ4JmtGxphUFR
oA9ItyCkW0isbEvfFbysWEjRYrFKZH9zII97T2RF9jvCc0hF2Iy4yuyIfEIcWAmN
/i+H51QqovAYg5PhrART+tDPrRc+woc47N/02rnUQyeR5W8OGcrIYaGQ12HCCdmz
K4+NG5T61kXbBvYaPJvOd3Y2CbUDCVzGZZl2fmaVFzBIftSySKXaj9L4xAFBz8UT
Od5SmFJFsK/wW2Kn/O5RNkSNOrOhacOh61QOSKAYJEcqmgozO7zxmrgGzbeO8sWV
1C2YnWyiUDOdKo+lqh86An4d4d81L+/wWJPskyY+I5IBe7gBk1+Up25yRmR5iXS3
z4alKGGRKcPDWg9NRM6dmGzhHPjRvXbW+LE+TWxej3Vq+47m4WECBa58zkhG7bjJ
x2hYCifPV3CQYk5FAE9cWTkKTlQOHOVeOr2q5Sivx+3i6iB8Qs2a1WRCjIzXyi5T
+5xKbX1GTIF/ZNJuX3+12XkX6wivzlNo8Dg0tvMHw6507XaawMT4mF8+vKLH76K8
wFx3Wy+HGz3olY7cFyr9TdMgIM2fU87MFNejVhAEWC/UApfLnDwj0L5V+3QRcoxV
8Vq1wwz57IlAqDpnpsi6opaknpFHy6gv4nADMXktDIq7piCi60NHxyJBaRqejLZR
ZLw6wN/WfML0FK8hNtKipmU9+t1GBO3EMZPT2u+Op9naxsbs9wP+pWuIhGD7apIW
lO0AmS52x30wyzQbzUVSeP/a65Hw+KGE0wyWpAIt0nHzQbBRRdqWKJx8l5IQ++N0
CZR8iwa5AO4OrziKnWEA7ZAQfYKnKgNQs6C5LBn3mKOJj4B909EqmzJkZVEGoccV
vMnR6A766Ml2vKE+ap+2RmPAUORiZlX6Jl75Q35RCm9kEmhiruf9c4Z0sUEUI3+l
JGGQXLUWAadMecQlrozD4hXwbCrPXpotDCdUSDvbuwiEYgvL4+J7j064NRS5BNx5
RjsiUafhF0Sq3ho8kXXFku88X6j0KQ1LURCDwiWRbOiCYpQ8+33uV8Nmr94yjTwd
Prcaje1GNK4hOxN6XU73wg0DHFbB5W5q3+4j4hHLLE8yU0oQCSSLRlp3qfiohY1k
/TKUglfsHSGKLELvo+HH6WZZeXS/4NP7sDhsJ4adBDnXfSXvwK7vzy5U8gtf6mZp
zQwr0wib9hpvTKxNx337uD2zm3aWdpgYoeai5zLjWqjQGgD5hs+qb9KJvOHfHvGt
0GLQAWAwVOtz0O1bC0nMG2dc/ZkgqLJiZn+nY93WjqlWFAEbAhZrtOgqjXLM3vmi
NWrqz0aXFsLwhLnHRkRV93AmllCMygYab2aOVfoCm6CXDdKu45/FjcwvEDQZWwRq
dtb85wxG9vEYy+t3AERZeMbRVGPc5EwYGL3Ni+H/m2NfTlKZx7HoYWjQFOE2LH0V
C7WZifLwauTU75JvszRdTlD8RxjUyVtNzZ+pIWB9DLodggjzFTEltsvKoMQyIP/b
M9VvxiruSbLpjmcZ2Kp48E08VKuFt1TGaVijUlEnRZahRpmPfKB5gV9qLfd/CzVu
uqt6clxfX+97Vl3u7YKkAxqlC5drc8BimodwsRRbPPTprIJ23u0LWUtM2DZq2aUA
sR+DfKxMMbsnmSvxr35l8DSWZpSKPk2/+WANtmfBUnmfmAcrHZolS2IMedcTAuxV
xwUjfvyTlEECpGtgiNnXOFmsBKf6TOva7+mMeqgzK91a6SZl5AwG3jCZSq5yV3es
EpHKgGgZTSYHBMQWaVMLfQhq1YOViefiLJbJlEt0pvLCT5eAwDn3TnuZDWyR9Ge+
8BGGYKhvEit6XsvTWIDYv6k29Ou1RIBM4IAT/F9ICkvDhc5pIVWtqAS1tiSs1LBe
oWPfgG6R7/P5yr8hcjutovPG+2z6pVRejKPXGgHpMy7DZLkdogAoI/yQQE5erX0P
qhtmtWBWbDPcurJJsMp2NfO5YsKVv8rOBf1rl1dmOn6R3WNgYnnEZhyCABjgk6KJ
t/eyKtrHlMXmwjuNGkg78wuW7opkNq/AiM+MjBOU0497vhQ+S/bNtYoS0gCFfib0
4tPL4+hHDbMhYM7VGgnBJW5QIx/mxVufoKNBtPvJVSZArKipOcyHRDpx88JFsMNf
srrvGvMWXY3U7uvJ0ZY3/UTLE69xVQMuuGM45ez37iN7UkkEIXC1TtqfqPy7wHG5
aDgmoBVVWsWeTbwoxkItdJWe1sKpinYmhtJK8nqeWydEGotquqpz034fwbJ7g3to
f64CtTNP0JzI8aXKFoXQBnRnji9SJrpqOE4PIlyyCf0DerS1tjC8n+OjJMLLCM7d
cH5Qi92XxXrB09cTBbMIxE1HSooc/9rdLjd1HttIGrEANIVnK/AIGOJ3KAE+bpC8
qc9lOzJv0XP5CX0FQLSkW+6hmSOABqVdYV4zYnY70CRRKkSjeIbjF9tSQhigeff3
Gx1txFeBCTyYpfGNv4N8uKjjudS0LHeCPPX4DAnDhYDgJjrW30vd54Az43cAxSen
e0/fkeZdqBF3EMaSCf7XnUAVLEqtnN15ETMqDIlimT2j86IMvYexSkXv+QccXxIS
kVpgFv+4zcMLevLcbruPEzYSPaGuNbDfLXW/1raRzntNv9/BATTN7pXEkrz+ugI0
7qIvMFethWWgfJ6Qu7IyyIXt4CGdsuAKeTWPyQTsukWXGQx1GYLaxfeDowV3gwTq
A4Ai5aay4LGqC19wjF2L3Bhw7uCGaIlBUULoAYWn++NbsJzqMikzSKLZAt6rqlRa
irRGhYu+hvSdTHyths6pSojal6D+blghzLvB4IFruNvXOn/SsnZaxiC1U0Y1Xfwo
qc92mxLv17AApBJL7UkkJPicbf0nO//2lQjQXKUh4Kqo3gHyvJjtHmkLc+XA0iH4
cU9RWA1qIvMlwtWBVq8qNJMMaSz3Q03a3VbQlO8mPhpA8yODd95w5GUQ+DsL+QNH
r84GlVW4PkGACGDkB1bF930MX4J68NY/M69+fTwdu1hldN7LRGNYQbXxwIoZ77Ra
M/z91zyMuIwTAjggliB3R6Ipl3FxKyaQZzW/BYB+OCN7sZ/Q6iOR87/cIEg62Bdd
hnZF5zmLTmxFSD+FWq0m2zMvJTe47/ljjaC1GlbwxHWCitu6U7SxbtQpNUXvZ6On
5ZCwSYSXwMz8VBFJlVEutrhwjgT99gzdMXOalnJXpvR+pR8lCz4qbjwmV/p8azJY
kbx2oc+K14E5LRS8aEy+1SauUPdtl3hPLTL+U0et85PcgajCgAadG+d+0BJhpJAo
MxdFALZTDQV8E+K2uN0208IW1wkFm7wUCdhj29RhxZQLFYRKk/ovFaLodTwDMzUk
c2yqcJZpstHtoZFU8vqrT7GLrm2fiCrtJr/hAMQ4kBlaTPRjBAmPFTy0bO8qAWKh
IJ/iyllqb3t2IzBZ/7x5XcE81X4CcV1DdHE4UNNLVoQSDhzDHE4XPbIKt4x+6eWJ
Nsw8x3HlJ8hxyB1yA/oPvIEknujus4LUpjGWCFnO+ms/c+SbSmEaWHv7Dkee7vIl
gx7ccGJox0hyihWFsellPf6rVixeL5lKvA/jE3kqi6xS/cq1Resp9IBQJyGx6Qx9
2ZvpqKROjjZfT2HxquqVZT8A/ZLSvW+uz9BRpR+cGZWq+Q7TfHBKhsApI0ERYrTP
RhSsomXVmccW2B0PMSmNAwYdh39ad9yY7R6dUCNuCeN4hVJRnr4MzAZIMgsM7AMl
mgwEA2prdLXgZsAHwWcFIgTpd8uUzg+oORB1+RZRpYqJ4+sbdZNXqkybmUflhJgR
cpeZqKVN1ceycenKucZs3WS1Num+Q3x7UqO+/t3Pe1Y1wZ9AtaU2Z24zUH2z/aTs
ir2nN3ceILGvdocn0bNMXPVui+UOizz3s3ZycgCiYVG9SxwYTiv8L2k/1sb4IMkU
1NF8AfGGKf9/40UkaPZa9mBNYFyfRMCcRm4vENi4NnOUbQHz/G0bO4lRJM2PFgis
nuhLpWYdWphxCd/Y6QsosHoq5DyjlrsMlOL3Uc15pjrYWyJR/0ZHIOtykUuC91Lw
0WQ9uAERyxAo3LBxOgbA1DoZJf54+pgv49uDdiESIj5nPPIeZvZPRJGEdAsTAPH0
qYcBfu6VkIUMHbk2l1vOa0ibx3y/UV6W0tLtuSAs/OABgdjLjST9zhAMJwPe49or
6pZvI5hE+XwPlj7U3qSysfC7tCD8CUfLBjfXWBNjmTvTE3r9YcM6I62UBgQ4Oq1M
eBFKp7WUz52neAFB7wSL7FNwfsQtOFv8jPMipqChwpbFMEYMtNwzsZ0MyEuLqwjM
nAFh+TDqamMvdP4QBbrCNEMgfh3XKOhRYKhdzmp/vaFgR16edfoAYWMyCcXBq1QU
M+sJmSofhtNV53PIJxmjDcBXQox21qMA+6cKmgqqJy/ZYVo0Immc3FlzLrvtUtCB
yO0+A/lSP85DNM3GiB/3PlLBUUHXVQGmN5P0ikA6xC+LijqmOPsVxzVe3WMIwFhO
1dYySC9oNvbc2ip+WtH1aInZ4rEiBVwXoxiD1ppKMDee0+ROieJX1g26wzfJc8kD
ZwOgddpxx2aCs5+TKJyT8uUbk1trID/dWunbPvisNQw35VC4t61yizVDuWjMyv6q
j+6zwBINq0tmDd5y2a/tdt3+7F1RQ5sXui6lvE53eHl8r9YrtR5ZSZHiv1YGpL68
ljp3J9Z1SZwKYjd+WnQK4XO0q2Bn+CVYkEpQ9fZEKuH0Eo/pn1BGy9X2XXmu9EcU
sisIAJju++m5o41mFBK99WObKnF1jOoy5wHoxbfrxUZJWzSPvjz1BhIkBqF7RKP1
2fZtjD8kop3CULB62OMttPpqh2lUXP+DPWsb1iVNPxuhOmY8zbctKw53M+GwG3Wx
crkRe4f1obHGJozPVogzwqmQ7RsPHJNhTm6OKfJUNXWq3AM9Ik6cOEGbTBZMH1K7
/6pvyf0owipOdrYWcaFub5pqaqcXXUhzWNGnrRZ1g9PYVJ1pvhSrTJyx7AEEGO/S
Ih7Q7jVADZaLN2yqDq325gGXgLdZ5+2GqA52dO5N4Ouh8EnxbKDsAA+84lO9oe2N
DcrIZjPvdMBt14Q5yknqDQQF63cMS1CHE6lMFKqoJaXXnIVObgv298g6uhCI/XlL
gBRoE1V1YbfP+aKSvUlWjD9c8qE2V75mfF6E7uSI4LbRjO/BfrlwvSQU3ZOkfQnZ
3rLTeL9UioT9rxcYdTfzdbTMJzQQiNtnKqrBlMvLmkH7uB4Q+M6z0YOnCbEroy7o
xuYi/6o4RYLjdmDWg+wL+tquNjf1toLNPczQ02Fac1R4QnRoQFpyQDO/jpSM90y6
d09nfySLWez798bZgRLP2ajo6QAHb42eUpUfNIGdY2dR28Q+JzDCSJEVMr9KBe0V
nx3fOveoTnUHFTmDxZurEOiKmPfwVMNg5VhdRLhFdSvJ5Vf+MTSTbO5fLsSeHTFK
t6jyhuYXXgvQ5+APxV/PycKBrEVNeikg//gZg8h5pExa0N1sZrSIX0pHhZAyOekf
wXfzQvlDGD0jVWdcZXL6HqG24wWoHU4FejRW174Ds8+tEH/aHFuys4oBwxLdljSD
m+I7Uy9eaInH+zRMzb4VVqRBRH+G1HvRre6QQZvYPd9Y7QaXUH5qeULTrY3MyCnG
1tXpPVbsG7qKtPY8MykV88s8LIbWlAwKnKLeGWw5RmZQmg5Sr/5m/GLWGdwBPoLH
6JYZZIua8hSWUhOUxSSCgrdNnn1jo+NWMGAvn10ORpx3aCJc2VOx3jZNcFoOj9kt
Tir9QztQHG2XyNf+rDEOdBCpQseOd7imGtKwAXpKcy9ZRUrvV68j16Yesdtf6nep
ka/nJPo1NFyVTz0FfdfQtD646+oi01OX3K0HzfJbecJRyyHmNnD0M/YiJkNj7+G7
/seXU6L/Djv9+eRe/86Co/1eC3y8kchNG6leoAB6E7LWWXjFCULwdRlM6OOKFHOz
hqs5eqw8LYh7R28oLTJO887rEo89MGJuHwg/zeC5bgJT+WpTKkHNax2maejAMOOY
qpaggcJ48fcnRFRCN91IQrNLWoRT05t4dqa7toj925rIHhm/xC8V8oGewSHYmv63
s8ca2Hh3yiDEcPwXQW/zCT2g0alDl7GE+g7xg2/NBWZz3XM0C5DxDmjPsObGoj+4
ONrJPFn5x1DKVQYkvYg0K+sXXy8cJl7kX+WipZL3sFBWes2TOD3I3Q8WEU3MTNA2
uEYHDyYYuB38n6ga4D/4LIR/tXPdV19nSw9GFwUx37oIJ6outiQvrJlpb9G0B+b2
3w0Q5N2tdP/IIZxhfLGWYe4s025fDQP8jvTE/xy4aKT9TJgQYgmpBJnD3OXT3o65
GwVWBE0z5SzwtGnG1xCgtCKHLJscp3o85JloxM3746KUOIv6sF4RJn6EYeWBU5/t
WaE3tU1v9ixFs95e+NNobUPVO9ykY9gTyNdWDVIFMf67S53Y3RssZLSJlUIfyLF6
/J4dkZMZHulF4Th0hMwJO1lXdcwEpm5h+ewYpgExZyhTypudsg9AwT4XsXQzw3Cf
YlWGkkWZM8lHqkaLpZ45m9qlGN8RBiOqN8+xqdBcNflufCYjczDoySMzd9WPYTg6
eghLkqwsehupVSYbYBYXdGTPyTx7f9t4+kBDY6SB/0zM5SbrYxqXWU94eH4b2GDT
gg/d/QJgb7Bgb7FX1lkMJLThEdEmqHlt3ziyt/h+/+MJL1kuQFSD3LdWN2MIaaO6
KbA+tSUiZRyx4RYGVKtQVDG4zkJtPkgoF4rcaLwHdu5SI8qjlh0DSpcOYZiw3m95
xeaQWJmeLEhRAZzk+PJrmjZ/YVjHUTzs/1yC/F+SmLt06IzGxbvPfwx/RtuQRPgR
M2tVjw+tsOQFmfjnIo3bqinwam5IANRsAsxqeWh9E7142/glBM5KDWDjr4Gdf4m7
taI7tvS5sWpiNa0Okoz9IG/T/+dsI589sW5LHFGCtSxG9XchV7MNrzLnHZGOxKIx
Wr0Yfw2oKQ1C0saDrU5EkPrwXA1jRQML9hRagwerZWR71YlLY+tChgUco7QBwZdY
0dsh4PuXCV5Tvsdgvj4BkxCIvbJhP4Za9UJvgMTHgoBQQ+m6F5E0GF/om9GZnB/p
oUcA7DVnrBsURhuRQU39aEZkbJiAA2VxdDpZjkdQJQA3r/F5K0JogrElSY7+a9F5
qo7GGG+x4KrMQxnyuWIyAnJ2zvm5wT2rJ6uyFTuEqgw/39mtB92sr4wC7lvQDhBh
6a87dOvIiB0cggzZFSw0mZjKJADSM4vQC7JU6/2sYVzmCfyQmIE7G1LEqhmG/ldW
WWDd9VqYz2pVZA2WPOuvOcUudCSRCy5XG/aW7CGEQgPwZcBWUPDP3r3byjmfGlFt
4h7haoptpLD0EV/7J7Uy7/cH3CmiivviEq8/KgVMMI9jFoTDyO6fxaZLZ/H3rs7R
tHg/tWjMKBH0ihFEHBOCEh1/i9dzLszuV742L8sVc++CudH4BVUwgve/N3Y4JPKT
lM05Zypqrir2C2Qvspe5gtVrtcPMHewc4E/DCceCsmuPxXMsZVTxwcx9R3VlxMm1
+3VS3ItSmObin7uDY+dCoSK+sHWeXEyJpSXSewUDoRUvp9Ba3RAu03SRqf1HGw/5
22sq8R+hl4IZu5ODAXQOjkDKSD8CBR4RYGH4oBYJ7A5t/jOaTzwP5IA7t2e6SGdd
9cb00KkVzdm3N1HQ1cEHus0E0rjEnXniQHVQhUjS38B4eYUJP/lO81yqVjxMSJLb
I/TzsoCRfsneS/SnfgC747QOdWYd/OA39Y6jZksOJGKn2pPCmjn0phLA8iaJM9Pu
aEoBbVvG286bIBBPq8WlEh/9NK+gFi7TR5qXwYstkIx1PHQpq7uuKy/NzBtffoOg
bARZcXW0e2k2CEJKpcZjY5UXp+479OV0hU7N89aFoHAVxjQbykXrOKWaDMqiHJr/
8A6BlrHskLfNzkqsdFaZo4SgxWcugUfkrhOxLHsa8tENRMey0GJkvYfMD6pEoG/+
oqDWhkR0W0ohPb/mrzc0/XuXzsA5zHDkRoFsVksB593GYjh3QgnNiLjcgM+40fcS
0m2+1Y3xPkFtXIjDYifaUtJokGbGDLFJbZy+OWfy++JcHNEKwR3sJZxNyfK6WMTC
eGblpiSfyPqhTMZFT5f9FEHm+IZZD30zn7EuxF/HANzvm1GG4IZpHbWobJkqp1jE
1++Aob0C3wN3FPPJi38Y0zt33L53SxAPC2NI6UNPiHylXoc+MH/nCkxUAgA80qg6
2hDa9sBAeOgxGwQEmPuPg8wep6VMUe85ppf72RxT6TWhod33Te8vQN2pNvalC6hz
Vcvm2L2AoS7dpZWyIAOthirgjE4/lDJeJ+sEYs1arqNRbQzKHI2hbQJ0M5LDzSBu
AaB9DZf3CkUW1gpjB7GJ7qc7f9O/1yNx497fs84jG4T86Kb7dmPDJa1kWIR5txBN
SNyc/NGEZH4QTxeb2PknwK+P3D0Q6FgSlzPKoJ20WN9ZMfZmjsHU1vSPBEMG3MTS
qOaieF1CIkgXsAQVW9OD16JSy9eqrzTwOMCt4WT4a/a4wY3oWl4MK+m64DIJ5F2+
eW8Wx+S3B10UmPfExbs7qgiM1gofAfmZ2GKyndykNokSnP9S3nrd9a1x30QgcDvr
quLQwp6URQwt8M1Sth1aeBA+kHbFQ+HXESZOwFx0rNxV9V0Uk8vAktnxs+N/syZn
LzZLawMyU4cph7MWW7d7LoZSj0tStTCfT7vRs0bxy1oTDDRABdr7oJcsqegm+IjO
exZ+vn7V4hkBNZpSDyu4eK4VOjhqEeNMCx7Ctm4xWPQk5w5axlJkDFlaDBmQIiRn
j2YX/YWZ85tKLQhX8z694jzl4vDq7p9VBk+0vmmRYJTzM5t3ztz+vdhtexa1B9yn
wIR/iiULwjkVOKFGqOEXTBbebZPxKTex8fLZxpAzBaKbvB+96qn4zMHF2Qffna3p
PnzW+cwM+Na8M+KHlHIrnlUrhIkUtO466OZIUQ3ZjFIUKrxtAC1lvbTN0sVmpjtQ
usxz4EgFTnaN3jioZumpYnZSHP/9g6d0Qc+sj27MzCVukqgX5f/s0aA+8c+0l6VN
5NAUJQVGlRBUMd58oBczFmDbLkEKZrVzNxqeRHwNurX0AoOB6VdbnzdQrmkUn8fU
yuyJ0PA/i28oPFzshED8c0CFnPmRBk2+bUvCyRMoOVilApGJc6FM/AAJQR0orFTZ
8kaWd4ydE+uD5RoqN0vF3+kbLQzaGQRfOs94N9RJRVGE0sQMVPv2VJSdFxa/6BJf
8ItO4p0kkzdmMeiZHslU3qFhmxpm4q+Xw477atMSp0Y4hpmYmMk695AFQIAsG2Bd
5LuqSTDSQwP5EOPaKotDLHKVb6URxhojsX69Dq/gRRHJtEFfnQ+aRGLRO2H9QXSp
XM5y5tj9wJEUf36vY7WAeweEiBtESZqWUkEQXUU2HUuJLjscKtWjZpRbbMI8wF3Z
9Ce/00coCLvX6MjrS2dnv9497kUXiuE43gOUseqnOpK/nczrnkQYTVOfFZuJOrZT
rCHAm6kaCGxhcvJHsgE70dPntqnJw96vG7csjAVsn4FbXwYDnz+aC/qd/a1uq+/S
Utl1jP1W9yibh+hFqpD2ZEwPd0JJ44HMVKq6JunNMHziF7TAIF+8LlhshFP68HoW
mkoaulArDRv6pPHhXF7ToINwl7UJ/tNH3hZ5Ux3m/44e+lskWOeSs2eekMh03sXG
kBckfgB0EWnqDHInoUyQlFlS5gSBFCrjs92HAWFuqO0GZiJuPMbgdRElLyn0oV+k
S+TYsx8VB+kYml3E4hovKMRFNPsErbsMNlFYZnPJZWMXGPY5gRwXSw+Ot2ur06LN
SNYHBetnygaWQqQ6FRzcj5WQASuXo5kwnMwL+aRg7lWDLT1S8kYODkSze0J5lxzX
e54zMrsBpfhCOdDoXHJjSXAw1yEBr6It2mdPS5x9GuwLm5RxDS935ymnm2dZyCVr
LZxVzmnuy8aedrlEgskYgViMFvKabYSHDw3BSt4DW9zrCe1lEHfUISD8+RgGg18w
Iq2pe1Vol7X8xwhzJU9sR7xEbjQmISMzViqCMCur/ny05VEQt74irEk1pV6NEp5c
4aGFtKhFrDNXx46hf+SqJYWT0GB98zEjdZlUw7yNfqLqIMdfcVpENgIEO3rF1rnf
sNPG6sAYjttBEtClQ/VA91lAeTymwRXVvHbf7dDSAgEo+PDGR+Bjex7viAIr1nro
eXELBC3KLRPmp8Nhiw1NI8PjCliXEPuCqxYSOw8tohVCwCPnHFrAzwC7J1xgpy7A
ZcJteDgdAXxszPhurUeTLc2+wzalsllg+4UtfwQrHxRY3NBXv8vL0/fPduhyodes
KXbwOUZgDD6BM7QsW/WMhjNMjRDLaCGm6oGg9bX8E0OHzsTicuhpK2/VNOP7Jn8H
gbKNcwcYqZ79U4bM8NA0C4pdQ+wT6xRtgWlCUl3jiq060zxoJL1X/LR48t1UMwB3
ilD/P60d4e0+dD3+7Tyt3vJnvLF9r/ItM02/3eCq1pH+diFVi5Ue9o5Dd+v0/VLy
XzU0d1BScd6mqfplMmuvOjChEqUR3NsLdgc0+vBAxLOT5Pj18QSCihlCea1rtGyC
eW9v8FNKK5hS0QnTU6YwfDqhgeTJVdWVOAXOy/SlWJP79f9MXlURbd52fmQnPL/6
0dGOvk6lpirqZcb2Su81Mz9Ee8LcD54GnJfB5Li2Guv2KIziNY3BkIYhf5RxTh7D
6fl6EDAJ3s2q7/TDdyx0PjFMilEaGUUvyTE3fri+gyRXDzzbCI3K+XRERFwNhohG
3lAQigil1hzh2eFjfuJm35Dg0ODncXPmD1CUz+e7ftCgIfgMQ8hadNPNKxvBJYvf
u2GcDcVwR7uJB5Dh31sraIvC4DBiwxceadDBLx0g3RbN6szS+SyvD/bQNRvlxnjF
PLNpAzWYoXpgRmTsqNiZeBD1vsKYrH/Y/F7DlwnjHc9+riXxl/vMVTpG15bSp8/Q
RrDuZNElIDH8OvF9xyd1RfdU3F2JChxZbbqXPzDJXoNRnhlhbeDQVmgAnq1YUuKL
mzu0eNlGzoxiV7mObxA3ddDl/okmOCr43MkklXXt3hB/f7ZmJRkJ7qpLiXQmpSyj
zbkAPnLhAxQYd7+i6W1qa6p7vam23LKhCwJL+uOlWCMjcp5lFB71x3rUEG4oz66b
EVHC6RKe/nTX5yFePSROAA2zG5dCPdvMMfXbIybvmejhmgLmfMFIOJpTqMT+AqfN
IS1HL+GPjqTNEYu3r3iY4Ci+vRlAD3irqMTv0AcMZZqEnoNoG/AVJ30/zX7muCyk
5IgPQ+3hcTeQ6XAqNldY4rZakKrpG1ctj2Ryi6UC4Ay4o5dJQV5tPTF2ooT5gHir
1LlzKAcH4PL2vCwpGfg17CVTmsEDQvYDQ56sTegjKEIzjwrNjdElgLYkGA7Nyvwn
6QqbgADQ/Lzz5LjsmNMYClh37CNwQ8GEH/L/zT4ag6Qy3bDm/Pblny9UGVdtEAd1
tDqnX/OhTce7CsFimbKiAlCusTY/Xw6HreRcJi+yKH9lJmg9gYD0AJCjTUFLTCcf
K79QuS6WCxXcQ0RLn2exWEQHqb4mzXITsYmEH1DXclrVC2a9XPWSSjB8Xh/PD4KB
IMQCOWQY6JoLh+ZTk25u1e9yDi/VXBEjU706UaLoz63cXhCS8PLaRIAeX10oUsdh
9I/GPh6E3teHtJUzVGSAwJVK+SD1cS6lV92K0f7l85D+To5ut5dqH8s+TmTK/cwX
/i12PA+saWoGy8xrtYU+3XD0ltGCNJgerS3kaUjPcs3uJn/NRX2JDAJWhp2r+hX3
Y1NF8hkU6NvK0NQyqDuTaxWg2ZvGGoEvTmJZtaOzeOD5+jpbGbWE2tPAJIZjw1mL
MqWugDsmK7IHnDl/yYFE6LDr5i28e0X9iorHRzcNZ7rIo+dcKDnyi1n08DxLGg1v
qqcDIX4kjglm8uO5w0wQqXBJICHX7xMGsQtzl1cnJ23/sdX95tANiP+1Qxp17c6a
7p5YvAkinO+Dl8FhIg3dl816/An22Hk/iiDysQ7T1blaUY8BZ5rGa79t8v/gjMHy
iJWDPGrmRBHVdYbwoldkdBH5nQwPPrW65/MrK6bE96yKuWLCTfwR094R4OdmgnG0
GZgNvQY+1HTPg6ST+vEEldbD5lJgUasPaIJlJX0GJ6rGxfQFpTGq6/O52jEzBb75
PbpoYZAQCP5oTbEgxOg9OR6rFndu1PtGjM+cBuNxWSEoJk4MoaP/LC3BfZqbUsZP
0AFypejv3uZSdqMlkB/AHkX0YNpYG1iTocwANv/UvKrixAEaDbblRv8g4A+FVHxl
KZD+kHodPUc59OlmT6/x0HDXGvkynw1mF55s1wXCLO0swJd5o9S7GB782nrJopVA
dN+k/UBdU7Xs1mym2qOjBmgbByxyADARh6DAiASfWzrnZJ92/Q7/BY/vcH9DMvsN
dObcrUWHQWOgeeLLSBqQlGSDOkDhL02GMm01suG8ZbugIB+zT5jDqFWoQ5eYCJaN
VgYU5G95bOOHnQIQxySLEj6oVmq5pJrcWUVpuKGbf5mnHz+RbYBTxCpQi6yQWU8u
2ILNg6tOT6P5QkJtQN3tth9QiK1AIkFMYMaROFmMzsT09lV2gQenKmyUGcxSFQr0
D/zFWVfDUldLAmJGexNmlOA0tapOWRdwwpeUkMDPT1RFRnxOuMdrX3qrUHCQkVNM
Vwfihk28X7OBJM5XHTCnq1aHTWmtWskNV0ZQkXZwo4TpN6/bIJNP73OSe4GOETDz
F8muSdmQSG3X9DP09DgaA/6fmZ9Yh5+4MT2ssPxFRTNYCAgbikS0RwttTUfZ2DEM
/vA052aAkBcHbIUh7GpB0PkAq4/jaHDvRGLY8VnV8mZ23xzd8sIPuqJ8yTA7u/bT
vS28cjdSwP5gkw5T9Zb/sMhOkHE7ZtyWNXDkJDYVt++JWOyVfmkdUYUlsT8Uecc9
pAzT0eO3+1b9VBDFWr/j4bY3JqrSsa/XF9zCgCHda0kJIImRhBcc/9mnycGrPx2l
3BwBYeGGMhtCgBjU5y+J6ZgrF5p9f2ej+KAwJnyN8lXlnX3/6o4Wl20r/1GWDsXE
kshQmwQ6+jFJR7UVJ78ZmiiSccKKQ1V0BkhdBmqN71YIdJYXL6p5wdAxDm1nawiO
LE+hqIl0PDdpbOygeB0dkz9fgFv5wsJNja5lQ14zdw3hc3rq2M8wDWZyvErwgZCc
7sE89TAhKJLDyUM3YQsgj1bJ+xNULm2wevARXC02QRiH3plbEwtlj6QJGEJh0xq9
FKRTOv4HzWvzuk0xfaC1KRlRsTF57SiE1Zjki/mRaNFSqEL+YbiMAVdZRp2iGWvi
AKd7gMNczGjsWrC5Ys/Jd3r4KTfs3yL5UmwM0+5qnzWhE4WO/eSMu3nfD6TBL+68
p9nc/7tuBmFTCK82UW0oGxbqLxWjGXNnAtxtXWeWr68M3qdMYhD6ie+dsBG+mO29
L1xoRJL/pochuaX96Z/KuwknbsBwojCHD8HwJxTVuhhkCoMjf9p6F36K63zfjeSY
bzm2w9xUXJmvKpfQEenP/YrmmYe2BocXccBA1p+g5KCyKldFJRNhqKhvQkYMVeru
VE6KrLfT1RHuLZ7lwp6dA+EzOE/Z1CsBrhCgLxU0eWGSyZgYGBaF29gijBzIcdG8
u4GoN6R8zGzOTjFp5cZpUFt77DbOQPRF+sfLBVs4I1L0CKvGb6s8UxMAH+pJfGKo
uUlvdoNEJ+WAO5oGGJpvObSfR2oKqAFElLjKfA/a4rRulaJT6vRqfcg5b8dcrM8x
MIKJ9kOvtR6CuJoCxfExWTQ2+PG8bGdkP6LNW2za7a6KJR1aT0fWjKBe+QMoRAro
afjkdPSkzJQeFp+1GSq276TRJQsz/XC5Rw3kSoeZzRhDSuceERHCD0GCzYbGnIap
eFCERPe03xFhM0b5gL7Ql7KO+Fx//WTIaSdNv/LMvjFgk8cjwG4rseNzLwaj/uiA
qSJXaVZgEMaSSDTa0tkE56GrxnarPoxBpTfbmlJ5tA0tb5+Noyz/npSqyPBqP4Ag
q82IBOgial0of/sF9+EUmSOvNYbEvSkRinsWMfp8E45kITenKYshrOxPWSB4fHIk
Enc/x4V9WcgIBmrap2QizuNwVZDxG7TuEdZEmJTOn2cNFM/F1KWJmJZatu9gIDfg
7lOvjmacR0xfz4SpWYNLH4fHq8Nz1Ncj9zbFQMzCbiki217nmkmMGKz19eK86t1a
XKmsHpFmf10ncVFKmmyD4ufVVQ7QP99nhc9c0UAAvzLlhz4hxXLUzVANLigSG1Xi
HdhrBXhDeIeCM25IznmJPMKl3G5vNzbSsV+FxsQO4f4GgZFgKBi1emu+LblfHgDI
de0JlEdxiJBsuGOGKXbgmTQmJEkJ9poOjCABUTGOehbHFG9vdSR72MIImJRP0naD
qrZcl3sOMxXVFoqafx2svi/R0/i3t0V1V8cVF6wNw6JY9srHbMdICIpAeX8k7/qU
wzbokliIRYQPs8GIqTM1wPkSUG03rlzhAFzFBCG/Oe8DdqtS5G0jMl7TmWWtGQ3b
txdq8XSshlo0k/kQNJpjp7//Kj+ISc/VpTG/u1BRJm8cdbeQw4QiokbSi4dh557H
exP/vVsbm4SCCnfPbt9TuH9IJV9A6Z/XVxsXbVf2dLTGWeOopMMS4ia9qyECBgJt
wHDYFuhpp7t5gDhLUX4cFERU8Q+1b7pj+SVGCM95TMNIs1tGxEt+oS/y2R9zJQhA
vCeC50WesptszFvpUhUgNvj0wQsuDfZqBmlm8d5xbKYsfc5RxfJHi2HF8nc4m+3N
Gm1PNyl+M9p+4b2BaAXiyV9bskbCCsTRDMa4RZbnvY6R7TGLvuwBtaJ7k58Ozs22
bkO4XpPfoW1LvKJpke5CjkdOSVdLjuWKByzNOnyhrfHdpIi5D7PCMvWX7az/+iie
pHlbFn8XkfVaTHUlssg4tUesyxXjuJWWlF3wrxt8+Bx1KOHpggZwLjOamVS/y68x
NMu+2zv3plCgc83XIZMqiLRh+ZNeAXEHzi2eNYO/ktiItGmQG1iSVpSr08m1Shb0
YeuMIceaVEKsm0FSC2CFsP+JCmZAntd/VNkFQsuGp09mUq1+ccDLVX5e484L0szg
piwpE2lZJlOlucEVf9soElxX9XBYhPWgNCqE4CGR2KNBhgpJhYE01v4f5H02S2Em
s/fffpcZIpY1FxTuEoFm/MrZZ9AP8wQa8eOU/tJ84jA/SWd/PHhb2GCUxPU7DLL4
lRrpDggwKjORuEIZsKuEtuXe6khs/CyCL+1c5Dx/KJeUnBPADTPsh9W2PH5sYIc1
RWofCToblxgS5DH9V1dNFXe59mucT6TnjcbK/Qi8CWf+jqA14pEQNskfOslkkcWm
bamBX2KXSqJUtZZvR0+sV4u6PpJmsaEEnrIQDv4VcF4aAvXFYxbKMfahB+sCl6t+
Ey4ce6FUzydkRtn6UqtFUoXD/AKg64f4zYu/8Y/sbBXhfWfRofu6OBlLBE8+F1bS
JuqN5WLwWXyujv9EnM3s6EfN53M0rkBmrrxBRzNcU70Eoa5bQetzmN4r0WL+hYeF
NthIooMu6TjNwBbNh7OhLl06AdvJlzZhqWULNYbaruC70w+Qcm08pktCy3xTKVR8
7spU1sPanfOJFgWOUIbJ0GeeI45gqdnmgN0MLB8on7piWHveaMQVJ2xSDUuKj++g
FmLfzfA7LaD0uoBM2+DYd+T9Sa3JVpQUQ98TUE9nT+yxm1FS+AnIhS8pYPD1EY8r
VJp4GoGZ5mVuqwEfCi7ZDLtdndFv4CLlk3oVsAC3ThO26qi8LQM4+7cgzr2xlDDH
OrgMXrGBAkI1h9wC3I3Qsceo3vWiQYCC2Q+dRz90ZpXaznM3x2Oy4eBcdPtPVOsC
poCr6nI3BvXMgwDv2WsESJBekf1HxL7VBnin6bFJbt62XvQnRnk8X+vMdHmtquJ+
uxKJRlzCsE0uOYOiejfx23ONl9ogdCOhzwvS880GmrX3FVz8I5uwgLmEq+DXFKWU
jBC10ydJXAUNSSKtq/VO7drDdcy3yMfU/mC4z9p2yDy577WgdOxLEWDUEzPvFXTC
HQJ6wDkCpad8drbDdQrs7RlVNbhEAs6gkglXdhr8QR5MGBRnisenu7tcgOn0+p+s
bygK2Hql5A+6fDm3phnsiC4JtM5N25ZuraH6wHSWy71MJXHJgIZXFdQ7oobAdziK
uxjIZI5X1N/pW2/AJ8dI0bHPUtXLnH+sFYj/WjNvoZHeQMv11M7vCxQl2fx5zd/V
On+DVjwUDSJzWdPJ5JZ/ahmorIG5tDDPuAFaHqz3HNcESbrnF9gjZvR8hIdhz+lE
13sC3vcr3/jqABQjR1L6hhRWDIC92d0QFJp7BP7l5fTuPGNObWJ1zMwcRyH3vXdQ
ZlRtZc1bOx1jsO9UhUcbFTkyL3QD8beoTNtm0yE32qEj5BzczpX7C5VnWHwa16+l
CiypLkhV5Pyic6Zc9I32/6uLW+i31fRItQpNO7BCGqnnZZIRmS+qb60Mx2uNZNbi
Os4+9qCR6RgkeA8095iCr4PMySjUKStGiCElpBF3VTn3cNQtIuZBFX4k6X8snT2t
+EOZ0k8dd+Pgu9Sex0KQPsMyxGKTlKSxfVV6LFZoSaOJYJUPmDND12saiL42sgFv
sXEeFjRsB3LMuxQn1yYtlobuMNWW9R4DAMo5/KhJJlFL93y7wbWO9Xvl8FAJpZpd
+B4gbTKikZr+jp5nxjoBq1mT19mlBCb5Vb/9WU3nwHpJPYjzZhKVTmo5eYviJ8/H
ktK13YHFkE8bOEInbkd77jQoJShzDEaU/kbRNcSlYnXnt0wLCpLr7N4doEBOb0vy
TwB/9pukpgmexA7z2tU9y8C/ASkmJaPbMmxMgxI7jrDrN+FeItJxrFBEA5E1x4I/
78akkLzj/1iVqYW+2/Nq/W90pNiy5ngRdJgef9SI5xjDf8DZ3kYkgoC42v2YaFne
wlooYpto7fiWwcvUxpmeqgkX+dY0snV+9foQsb1iMvenk2fVIyv1GT1mwu7kaPcq
0ETp05ZxKZUX06w2T5Rj7hKJ0SHaElXeGSaH8FE0/LEny0TL2Eby8eZBtrEqZtuf
ljt8YSdv1mizmWaxCb1+PU8fFngprQgvcho05i4lnU8rbtRpPBWtiO3TDhNCJQ+O
IWVxepICEqs5q/AF/ETEcDWgjmmn1EyX3g3qAQt2iMgzR+GJOtZEc5VGa42HPV6Z
/KsbPhB/1J2JWaJq25wykNPvqLG3GMqivhlvDa3VY6YEBNXRcGsdy5Epkxeyqu3l
hSuUNZvm710c34EvcDKOKK7r7mjan19tF9dKRwJtAnTFrBLgbP1OUWGz572zvAxP
ACcO0AwE5slpc6l4tWG7pSTfAaiAvmv3KtTQ3ev/kFfvlMyBvw2seavnwasbUs2f
ZTEulNDqHsDt+wwDRaqnRDsV80LUyxlRMx1vVcR9BReu5HbkaF133x0Cez0j0LoV
X+zkPLvvo8xnnWtDTtByIqW+Cd1LZ9g8ne8xemU2Ef9rdEzwdqArxNcbTzksxvqi
2ShwGMiQFIkliOEVI/ZUdOk6bE+X1bNpC5+37klMTQ3qqgNQestQPa4/FsPJlou2
J38/IapMVmJwmGr6jxC04ZKDY/5RS2R50arQ8oeRljiD7ctM9/t2gnWaUOEccVD4
Z6s2YD67F3KOBp4j8F/HFRR4ngAu5ptPTgbj5b3U2J6khCy5sDu5BoMbTqK++mD5
QMx454UyRlHH50omXDFaWXZv/AaNPkmk6rUA7lxL2MyK8UwWz9jrZ2xlAeCNwN0x
toFy+D00AFl/xWXKyqW+9mDURVYTCGeFQ90Hs18szg3HY64QTZC8qG0eLtoQLnp6
VIEiDU15x4E6oZc3Rcwg95RSvOzGKQvJ2CH+TMmxOtSP6FBKZ6OlryOC2FCzmAgJ
6uAfcwOF6RO/laUB2xsJUs56SVE5dC84lfLbDTkTmAzb+D1JxnNvj9q5OpucT4YY
dKiywl72ZLWAwIf2hAzPTJZ6VApzZbGxJZ4Oa7aNDVEo9B5xjRiOxvFWit4LV8Bc
k/YfyrWS9CWVQuTr1yGNLc9Hgg2tiRxhrQdWStIEbQMsq/5YylphyRORXAW0Wuvf
vs6ppuvVI+F+2pJ+QoXwl0lmbYTeHvLhT4C3AEyE+vwQjbGUCtVdOB3YwwDGNIQr
CMw4+TIRuqROFYqiZZOGJJd9GYrN2TRXyAyxuZs19fOBETg3e4VOvqJs6ui5SQPD
TEg4T/yq1sbdGLZcEE+4jEJO40D7vJsK5y3SZO1TDijac4DBl/Wcf3BxD2vMRgzT
EfgIr7kHB+SJrzC+5vWr/kOLV4jPZYgUBRR/KeAPwLuATS09CXo6+O89PDoyZjez
9S6W7B+cbs86/yzli7iJDFvN7IA3dui9mWL2nf6b9DI74Ls07PPVVc4qwEXqqqU2
1h0lBOp/Xcs7tqKRszVEa4YPYwgcV5X00ihqAzZXvpv7c3iOsycDcqP+1+KX5s9O
jfSaog+0dsUuCMf5JuBeUrtRS7dxDKGpnIR2d3GEyapCQIl62NCgcoeeStlvQbzT
kDvbJ5Byvh6C8gUr99L6qWGmajyXyvDzQIdR8/Z1n3GMGk6GMySScDuLdvcZAdxz
PI8yhsbVBpuRKUWHMGQ1edz8KjJfvgx/Z53ZRLsEzuwGwew/GkzSDwgAmjtdEop0
ymwaU1txImhfAqi3LfTububHe1vbngXfV2tTxOryfvDgg6/6ir0+D/hsyM1/X3q3
f9r4VzQBi5VqOso3nSrtQtOzcostfGKuYpKIhvaOZh8vq5GihPUhz0o9TE5IaV2I
ZkM3xC3aOdL2etvc0cxrJcZp9eImJGyPc0NHm/g5SVBj7Ts/b64wLTxeJSHkf/e0
Vk5O33kIgu84LW04URMna5yw1Ymksu/nNkUrguEMg0QAR+dyUEZ8WqvEZVHAsztU
zP8S8B3fL+z0eg7J4DSGrlXDUVYRrjrTkFQPLFzH578esdC5CPiikapbKRhTX1li
+YzZiSRaNlbv0enndi0swO/0bm2Vo8n2qmvu5d7oG7/5Lzrwmbl2/nHevpIBOalB
pR/Xm7CugKUF85CmCLu9x0ByWstmizX6mFlBQrvhUd+e5kbhO2BpR+o1e3xVdZz+
MwL58xUXw5X1HqOn9M5GXs4C8HXViaUO/O3vdHANCWxLo/uJDn7obUmRH5dLVfub
qiIWQAAoeVB/KkKsinYa2PRW690y5//YFEUmzRaLbS093091X4mfzQA9N4jeghU5
7RfV1jvVMXeRDDuGK9V+OInDCM0Aj6URPo4wt2fIPItgRDx1l3SQqMGg4JV8kGO+
ENnP62+wQQTwWncyq11hO/dVG7kevw4a6Z/x2w295Wqh43xYuTygpACPfy0MX09v
y99NfCJXqtO+h4QGF737NiXySh8ldiFaphPHDC28OLj6ZnmWtXxrJ/Dz0GNVL4Qa
SmnIPQaVVyTLH+dc/bMU2dL8gmIAU35rm+lTUtJcRJsTfqhWxO9Rv8VLHqep5NlG
cLFoNg02E10Ct2fPe0UaCIyoMRJQrs4ZvG+LweYO+vCx/CED73GBPEToUmO+NnAb
tM4HAcK6FRianMFnJ2acKZkECe+tbVyHE3Zm8MZrWtS1YPuxklk29S86cW4UrdzG
Z7qTlwkib/2pSgyw14gbVnQyy0W9Pp80TCEp1ZYyLPjFxLV+NNkd0Hjb+T+29BKc
/C5XIP73lRu5svft+fegchwBDG+8foXVYv1c604fVroyEbb+i3dU/5+fPn9P5zO8
F18IBTesTmgLEC8z8ZhffSwuv7l0soU326705YebN70ETuGJOtETIlLAFIi+h0bC
g9EB8ntkJFaC49uFL2zql1uceNQymg6TO3ogF6iM51LusJGkqmV1yuSBYYgLLDgK
NiMko+ag7U8n9k56RKe9dA8PJI2P5MldZxa9bApvqD221zRgF+UamMbgFPzEGJQJ
padbypB692DR3qruwDmEkA9WVVNqQMjGQWdy9ltrLf2+tmYVhtil4G/Y0rDF95id
4XM/t3/jLENw2AehsKSinK4Fw7Sju5Nxv5XozgfrXmJZQn380Hka7Ylr5N61njHU
cgI09GvtDt3R4NltwIyBL5Kj0vE1U7FU6YgPHwu8nvS1ls3vEzJyksPSA00LDFaw
JpO+zzVcSDr/74DBBSOYrc8Uf2W86HQNEQbZKk9LVl51qAVCNk9rwZdYvODf9lpv
W55CcRY3dTgCKICGNL1tvBuX0ejnG0VJkyYZDqQxlUsVF5uB1UPifFVwMeNvI8us
NWymKYLKBxRuH39qBqjT0k6tOvDWhb02oF5hrkw5Hhr+LTrZEZFYMRgMhUNwyiJ1
qCNWEl0T6bmlGOIhQi7d2JEyx5MEEMzysWNY/YhBLtoFPi4aWvITDq3g7y4P3hqa
od4IHVN1XhaHGYNhLVXOpseu0dGDyXG3J8clkKKWRId0Nsvfiq0z15YW5XuiRntt
dmQBOI5Vp6JpZO2WvTLZ86loCR1bnne1KPyFoiTav2d+pSxhiq8eUDD5//3m+QbZ
jJvs4VZxpQqmYpri4jBai5X+f1SVzRkRhJ+DsUTng53HKBOgy6YmQRwh/xqUC8mz
miqJFUL2gGnEzYScdiOa2YdPfpDf8/lLur5CHIR66Av0cjhNkfEe06lSkRYm6zB2
36PNdVK2Km1dLtiYfXGZ0iaIL8MhF/TueoOHhTwU1CPr1MRVALyILD2g5HMJyE2X
hlWNpRvn2f0dj0RWN8u44sqSFrPOirA36qjvihv2eemMNeM+cV9oYnKuQuQM8+ZS
lPc2ZdUBpPAH895Ktffoys5tG9gFXkhmBAv2OcUVIBPmyvm8iQ6zBrAw5aK5eCEr
Y+n2YWRbK0nwSPLZ18LS2JFH3vpLODCfhxwPwyxS8pPukMRppJrXnTcfFCt2xkrU
5UIavfOGHLXdaOFgfcYhmvPFrujqNAfRgj0E5+bsRLNQPs+zZ6ljKaHNWXRDv+/q
uJ4SODA558mqChxtthkWQdqOPv2szxnz4EGHr31MHWxA2DpMrMYqlDxU1mWiAkbm
U4z561NJcOaVDJom1UQbIKk+wrOvcGw+ozVejzJGOxyY1baq8Qi6LcHSm52BwndT
fdiddGkxKsny7Knn7y5SQJXFV9RUGYMcZgnbxiFyRmHXQXvOettUTpWy6jXix5Xn
IOvXlS6rZMk5chIbBSo7Z8bQOoJIiR2wxIoOMPLW8rQ3cbhKv5Ur1tCQcLf4jcua
JaoAf5iO4aXRFbUUe5mtEPDOgjFqhpNGxaKfXjFZpjCXUlQFqTtj6N7cItj7tGwt
Ox1REfv5riwJ0CkJu+PMpN43AlPMbFheEyDuhvAFFgYmI96DZbDI+nIG015ehRIr
q+5u7vljfkZq2xHtEK/bH2u9vbGdPJe1g7Gv0WcHDW7fvgBWRJVmT4Ptdq19Ho6V
cyK9gw5wgCBHLlfsDNPUc+OFfg3YYXZyiwhmEp16O9qD7nJoZfY8+7J5318C5Kht
M1Uy6SdvEgqVPUJu6gmW6odFjigPjo1555RI/cvO/cA/2KH6Vrr6sa2Q4ohyz+nI
WRPPwd9NiQIAA4kl9kNZqRpJdOdzumhkdl9loSo0zemXPwQ05hIWE5FfAs93IP0Z
sqCof8VR8l3Y+yT8jgALHS+vL2735QI+SDucn+LcXp4Yq435MgXT2Jzze44oj2QF
1BYhzv4yXxYIg+lz4VP5DDqnEvLRRMro2YJXMaEs/DN4j5NZOP1hJneXqyeWxrDO
p3x1VMu712yskfu4hbww3LEGIK/5BOFnz2qLsb/TfhhXNoOIzjzlxK0q8WnR4FYc
3OaazbPip8IMk468XItq16wVlCeYE1VQ7ha4k3OsCoHi2xuZcwmuvudbTOxwcc+n
zH0tN2pVDJCTMxw5ZcWTDR6ew0PVyLQopTw/lkVHNDnkFhqNVcO5Hvq/vnfunXq/
7Iyk/EbinMCRtFQvIGnD3Gf3bFJeHvlDhS2u4L4phZhAwHpBM6jg/ianY2cvnH8t
z2FTNXXvQKl6nWNke/369snYLFuvk/J/lDh8HbVtGlmj2WcqvtPVZELPap0znGB5
zrB4cdwC9/KPiq+cYqffUbKGSbJkGhFqyOrKPfQCAxG8c675FMSEnl/ueyPCh3Qz
rKG0dIFuhcd5TrOqAs1mClXBOIvoGBUvZyz7Dkvad5fXlYAxvVIfhkcey882JQxJ
lArsb9lDVH4bXAwDl0FpwMHDJ2x7993nEzSdQqVLFx35FBzSwvK8iNgd9yxOZbVI
zseq/nnQIyBokfYRSJp24CY4WjOX92TEwYvA6x+uSfcwd8nwaZnIyi6B6O9dfPnD
dQJpIjuLYjUpLAG09ij1BgEtsAiYjB23z6BhWjwWugPI98csfHPd+aio1w93jXND
KOIDwHzehTnFelI/pB28paLLOA0Mu6APeUE5047nMCJsP3MoyiBQq4mTiYnJK4L4
i5K6r52uFhAE6YO7aqwNUi0QcjpCJx2veffqfjZbCWVk4OjXDZAeaBvcrxg4zaFR
TLkiqWPRaYZqtUfWW+j6mAc1KvV3N9NME6jNiJbuTZbPuB+GoMlfIlVToS/aNPpf
De0g0od4xxBjTkoV6jkXFUIZgpQaFrX2XRDzy4hmKxfcy9cTHhpjw7iHJkn9Ioha
dLgSdaKxF6rmeoFS3OvU+Tsx23yxmgYCHbjrNv3je+ZKH2dJUp24dx0+suFfmjfd
iqr3cHOUHCN6sy6NpmkWY73smm08Atyni8/GNi35WAXJQmr44PEemMO/qobso2IM
ltYkIW/pMyMb+231nQ7wGSq4uHEsyypDxik/5ogDf0lHThwG89nn3js9GEbV1dKE
veO1ob+vi5RIoWK5GkHI4VCRL8VyLVPoaB25dizxHkM8FYzzpKtUwGSI0b9n81wV
H5sDBLsk3XnAECXNwpxStyp25nfbZRD3kMgCk9cwPSKHbBWgedQULQQ2ZuLxHKs6
EmxPTpWa69Eh0kyDc1VZcDmTbYU42MW3YNDXzmSzUadU3iZSDTSNpb85HROk4QUD
uwSx+MVvtTLWyXwrfoOhqNIkIZkN5mYNl7KPOMbN2EqEzK1KpgOxJ33tZlrfcw2v
phnmMrt8nDQMjMbGHBCe1Pbd0644LYxlFwm+zSK5hYZuI1Gtts/S9bpE2eu+wY8R
6KUUZ9eeUpGyLf2jZ4gLSvQqCBu/3GUf0GkcgRgxsLlFUMibn4itHBflu4suHN6n
ViKdziChBTpyK+TSgsiOH29zR/tplKc8jN42d6iWpUiBY/5egDqbQGcVUq62HnI5
V9/ALgivP8vzHtG8Qwr6CMjUFjYRo0MSnf3wWRNzUlS/GYN0URsxaHLVdkgwfChi
razcxyDFTO1DSMaBuGkUuwTqliJxpUAwTQa3sodKFvgciVwFHYfM09JXG+z4qzCu
e/DBPCYUf+txUVw2irA+IXHESbqXCNX6AYrdt+EXO4giXgWd3gwaGsqJAE8Qi15o
QvVztEfi8m4dg1fBa4b3Dd9Jo8oIVVxNLp/ptmCiSo2MhxhVcL5JCBsQjU8szbqI
loe7EOhvaP/zD4+ZrNMf8SPYeSG08YW8lE1M6RBroYSJf6KwAo1GDWUg1gc04mLg
IlYDM8doNzXqrrXDZijhfsxlUuY7X695IDwigJ8oe0Ouula6OPCGOaQExuxVqwd3
6jqbGWsCZrAXq36KR+g5IL4OllDO7FK6laVJy5kxsUFPN8sAI4hOLFSZS8dC3t0+
0U5T1tDLQfjAYzYINaL8uRJdG0JD5EkSshlnK6cc+soqqt/e/DAep0Tg0vI+f6We
RXTIWCcwL4vvuWCdJ+HYh9rR3RNtJPxDels0i9ODLIm5O3WaRfb104eGfVbiKpPi
goe36OKzQ40CtObXCisqnbuRL5kDggtR83kNgdWX4dIgFUNYJcSil+cOdvg+ZO8l
x7jtvVuj6RETyc7y44xmvChW+Wp5zdpvqKXT5CWTRvlpK0tja6kVe3A307omJgCf
OCGlVI6s5B4Fs0m0L4l0zmXlU9LxRL5Ho5KZAJVqIuCPAmJPMsjSF/EfkQza4uQj
0j2ZRPZU54Ie18iEdS+gQ6ciCUXilqtGCEzNvW8nEJMhqeB4NXDSAQT1ukb6m2yd
kwF95N5swD5Rb9d+2SxNaW9mhwS2dugxLafoOraA4nISLdWNeS4gOXU7p90CDGx2
wOZa41JT/4yQrHeuN1j5MKoKmTv1/DDihf4mD4o0DrBIiHRBTosZQyQiYKeNdEDm
afyzjkFp4JQo+U4isl19H8BsdHRsMrTwwZ0CTmfRao7kdWrFzjz1o9yq+0NPKWcM
iX0msMkRv8TvIdnzwzEBjt6nN71sELdT7t0sYv8JNvuLbnkCNEkmfiaV+4WluWGd
r0FTq84pVxLY/R06ItkzGKn10uzxO9VyJYiX7AHl2kJWiz22OELpF8/dkHtfrWtb
Pu629MahyoTxilGdaoYrVbqRKEzX0BGO1N7pMW877Yr+9fyv1ZwaaYf5CYgfBh0L
wZGWoaTRc4FWCFZi6fwpBtueTF/hwzoIN0y2wrRPqcuOxjZZSvY0hyrmYVPjjzmE
eJmZBkj1shy8dyksWvFdfmMBvVvfxaiZi41AYLR9ynQOUOf806T3A5gSx1IOHoA7
1DJv9/frQkMsz6OaiWd/aK22u1X5NF6j6jkuSvfX8j9I9fxYERGtlXFXjbJ3buxh
iZf91ZfLHvFxOZRK/ZRqlWMYjQ+V6Rm9fQJwXdoUyhAz8ggGlZG+pcrwpO1yGYrC
yAuiDr9gxrr36xkpdxiLrywj7elONY9oiXx2W2fqsDZkkpj9MEzZHxUnCACH5pRs
wgiqvVBcKWu4sWdAiM5hL2fMBK6Qr1Manp2EnLgJXksyNaBUcwSXVA2tcj6ysyIe
J6GCsx59QR9VbwDyJxXubSpCIg3BCx2SYA2zjmB1O1TF9fRNC1mPT2kOy9eGdmNh
ba7wyWHhFZwGFvoLBV30IyykKpwuf895KV95BLtCwNEgQ/rz+i2gnxXkyHjV2gRT
2rPDy9IPvrQKNuPmHjpo4yRRLcbGZ3BBdjWocTVrffqOzMHoQoIAU+VjW0ss/g+b
dCRrZIOc/8NrEoPXCkDYmg7YgNc+k8Ss5DZsSgqaNDd8cojSpa9i4GyGyuW9aGIS
JxBGTYxiyub9KoCt8WZIJdCigZUFuvT/QeCfPeFqGbN7Uw3J0h/xwlNiguqq0/Ne
QdccD7LhCLf7EL8PLf+DbQH3m8F5CxExfUxzOAtHb9x+uDMLrsAQJ8gemi7tApFJ
qzKq0capa2SpSh5pSbmxnnZ5Bl/BUYVvjeCvdKNo58KM31A9DKEea7cX/0AfSZ9D
NcjK0yYtkeLKEWWxkbuU13Lvm7Pem7dCKc0/RhbPHvV8Rk/ROOoGjVBXGnErqHqW
xL2KbaF2BNkWzcNs35k4Bbg1DKBXkccrme4eufvGTk6pMbWN/8VvtMjZjqF5jH5P
X5j4a29h3ces9NIDaD3k1Vl12ADze9waBNzBuYQiuAkwvLR3IlKj2nYRYgah7H5y
kOwASx5xBs31SgflK/4niTC7rt/XjQZelR49DpeF9zWs5uXtB6aimhQEjCoO7xMY
U1NhD7K2eb3DYazbHQy2EqH0aa1IAgmfTb3xggjxSZOAiE/Xsre1A1kpFRGgYZLH
qFTtakzm0nsh/RAhT0NBjXKLkvtQSbFQX0eqTajyxZOMW18tnFYMB1H9xz3RYou8
LFLJq/RCb7iSO0Ot1epzT6JkuHxbXSBCIruoC4o7GhWE27d/hYnT9PiqjBfjZrhw
ieHWHJZSMpflRAkL/kHqRn1LkfAjeb8Ii87I4fxfBwl0zWYWuKfxMczhBV/xo7AZ
VYYndkn0fhs+TKRhBTSI5Q2rZTYuoH3biN3s5rNh1mXNr6Q5KDAza9IUX27CERvO
YcPZ8j96hFSRcWR3jpgq5UUioax9o+lUYlqOBsvm6kLdZRF080INNn3C6CSp17nL
Rm6dlWxvmKnbCYfdVfg+mCVMXqR72xkkEC9uQ0kunAclwgdvY9PrOvE80y9nezGN
Ez3OPCm3vSdve/s4gUqhGeHMnjDdbZ81YPYls7m1/e+TyQsbCe22EJ+JxI0tKuVO
GDEnYAibCrQwtuTpvv0Bzc9A3Cey9bs/NmCotnGna4PIIOBEgCpDY97RGXdh+bsW
VW6q9AcnkIIt55yODdxdoqyTThwgNehFUuh5Aaqpya36dQ0xpki+YssJ3Ke9/i2x
JLxVBbe6e8u8rE1yZr3hv1j5jzyBAVa9aGOo3BANj6Q8GlNu8olWMtSBV8OJDZBg
v1vm2DfTYcB+E5LndkJDkA8GhAvcQcjAMRxFDhlhdPje6/q1IIJ9hpeA036LHzCI
7/gG4itMi8HDPGeWWZBOURs3BOGGMbO0jxBP3sgRuwRMfbMLLakAbA53ucYvVMW/
7GMq0uYskRC+vJcfDOE1zBuPdb/g9s6n8IihnvtuK5AqGTemmUm5+wIleEtQKpi4
C12ihjBWGixHAcVsNY4HTts50yiQd9zFf0AOf5kX9A1jjYWzFZY8uz4Vg8DBXKB4
FD+FJorlDNwNcy4PIAtXBcjHNDb0zPi++EF+ANosX0vdfcXGfLtAjrF4neGW58JQ
284w09xKzIDal9Y1ocPps2jFYjEHC9X6VWr1FgjYbdvtTNCDwUGbbpslfOP5ewVh
y7fv1lvWHJYyvGgrOcBApM7yMj/2FEToSGHHiuHmrQ/N05kr8Pr0flRX0WYqjxbv
p9f56LnKs6MP1Hc5ifZQ9jv01HUtpS20HMqNNGMtHMQgzmZsvGJcVuRxc9P7uk1u
3SEUME/uJQ9UpgMnVwrV3kByk04x7h9846NGN4A4hi9WVXDeEAxAKyZ5oUTFpu9Z
c6rX7uXPBGRUwfheANi++cubTiLDrJeDh1QhtPJHJ+RD469k9aI+PAOXT4XoFRWB
dHVAByaux3RoiHF1aCuGZEq+NmrsxZJDjOmbvl5UeS3T/eqwuMv8QCxdneG9E77X
xDDizKJ4cC33MsSJ2sqbBqMUosc0D+dkArt/89miZODAfcoB8aGFl0o39Udr+bwc
AjvQsG9awP60p/eI34gM5a79oekCV4yG0Yq9uzNetJRS6+YWP6PLHz1ikSibatVO
Gxx4EcqfDX550NAyhkH8vZgDyE3oEPLWnfbmBK3SVCmD8bYvFQKq190WCPkAy6ub
wWSZ5aCbWLoou/IlERatDXSGBiz6DhdNhGz6/IWKDsBwfs77mmVsOGmTArptH23C
UWgSM3kRvWGgLovyE+yPZ/3uj7QUQ+igzCY7T/uE4Gd7NKZYxVfzxhs6YhDo6s+m
uMYGojvTdA33NlxzZ3X5PjtN9oQxcQdlAft/t0vNHfGHJBfQGm/0oBIlWQXGSqO/
ZbFSyJ+BQf3Xl0bn+2dhlVvQpaWLrYtb3DaanJO0Q189k0IokfjNI92abFKzpZNo
eC7B29qvdwpMKxSsLb22p0BGEYjaUHc5kfhI4pi53y5anUxFBMnvBTGrM2pRWiRp
dCKX1615vvVspKhtH7qHJeXk7KJsi0KwBd/2V12m6ivXqRocgNYVbijrM+79pFmO
xeIrzuk6X4U0UCyuT2d9VhqJdJVkYvqUeKnnV2iFqn79eqHhnp4nPbSTYIc49SQu
g30nU2Zk4lioZxgI+MP4CGtLPMxG/H1l+FNf+MXLJzSzLkvPUBoOBgM0G1l5xI6b
yGJhmdIjYVJ6rlRUvAnSZkVv1F2B5y9ocz+mj+sns2p2+sb13jp6lpHFlG+/3ZNJ
IF2AyWwpYl0oas87l/iKH3DE2yEaYcooRvSrNuaC8VIohvULK5r4wXXoDtt0h4Aq
DvEpgPaoOLLm3irLxSaI9cr3Ms9xFFg4mWAZ9AN73UqqiTJNje6peqXPtd5H4wiO
/hFPbxCxEbRwGNA4cm0R2pMvjkhadTolY2/HHrWWNmqhVCt1zQfMDIXV5PXyuYd6
u2fCoPel10xYpQeGHnFvbjl2TwM1/oXF0es4qzQ0vUkfqPrcLAPT2giuVH59hwse
TdI4ZVgZA742/ptHldEcEp6y1V/laslo/UhiFwFUzzdSJDnEn7Lio+SiRjt91IxO
Rb6HWK2zpD7/kMt5xJD89o6IN33oEntuTwlwOKmnArQku6e494FuwGM8LQzDnfYD
iDJP4flqCW+TRi04LrV/Aib7QRlCxnl2b3DATunyj9/OxPfnnW2iWP++ycQSaLZh
UqlRxEiMag9I5dQ5mN/FQe8BnnLM31cKiXtGg4k61ijCmUEslbD/VaN4fuZc5Ghc
kaFzJPU6B5VlDCjLn2a9m0X+aacg8zg5nkPyD/SRWlbdXlSxr0cI1iuc+UV6HZyY
azWuHQBKx/w91qZY3ifbwNIJnQvW5zcYAUDmVjZPWLsDQYlIPJIU0BFKAAXq+l0T
oHFSwlm1dL5na66dAhmPqBa43XRUft1+C/APjqj3EnaB89m/m1wsOcnjR9NNw43D
Jfd70P6jDTAghLfMDoflxB5koROWk9nGV9bFVXaszKXwnI9yYR6x1Y+p+W49fmQZ
JBvq+CrasaDHqI7OUxtqxE5lX7iAYUNWmRLn6ZL3s8ndI2eAWjgSoPhqK43CgLRi
eFt+8ZXDKmnTqvqSFfdtRJqpi/fuZzNUgcPCUgN+dzCW220XJuyO+z6/0zWMHald
FHvt6AXhiZToq/LDo/2mLsxA20ykCQsgXafCUAlcKPc7LxlqJdS1Qi8niYVR9nqm
e2y/d1ZOiMMaLuwPcEhUXJEg0zFos7Ogc2+Tuc/AEPdb3eomO4o5zeO8JbmEikNf
R18Hgx18Hks+TuX4TgftWuK5uAMJ7CIGvU7jJR7MT3SkBoD16zYVsMNEoFneszBz
BP0HvjYJbJZ9kLsjI+n+9uf0DfyrSnf08894xCdRhFvz2kLoi21Cvn75PtGYd0/s
2/kJi63ujVgTkZZalnyQ1/3MKThfsM6qkMN57RDRzD8eOkuGKI2clKXtJtL3ueYl
ubYEhkD8s5Ey7GsqeIpyaqo83SCkWEDQG5kmV6CYXTLT92yje/yZPp+AD+4voVEW
zRgAPEawZII/tQD+svzkskFnqDskW50ErS12d3eBqH024lqTGSVZsuhkHbSBEHLG
9M4qPy89+qHKhgx2InBSPy/n1QVz1GSaLdoK/G8vlIwQo/q6vqRtf7mhyCIjdYrk
q2XNOLwMkDOuiATnvXfzjS5bibY+ZCOnjaKw13EvqE7YCvuZxTWRaCamW68IaL0J
5MJdh4sGgN+rHdKDAwFuMNvpMCv4m2kiP7uRMW0Fmg4VAZpDgw6pUc3gbVBVYS7N
89XYnAx38abX0ztKiCw8ICXcyKKOYpnFvnpuKBuW7CWz0Q/Bn9H6TxCSrTIWgPwi
E460b2m1/LUS9MFdSrfMdTa5i9OetEFlWv7QLn7HrT11MgLlXWjaHLIKVKOaLotA
GRIL3zP2mV/ymcnD7mccgZxsQLj4glmMxGFmhKtGGmtf0k/m+dwO6igFIikXGdpp
S0FBGkhpkUHR4rAAy+/zphyFffWYAU3VxTUwMW8z6suLaW39XrCALCVnRqABmWEF
m9oQr2uPK7VKWuS8XJjk4GnCxz0GKZLgH20TIl6PIMb8hutMIJj+BRJdJkP4jl6Y
n/slNULsgoiiBSxFfKGLelNl6tpA6rO2uuPtDO5WM2b1ybbYk9no3K1EmIRYKVfU
iX5bkoHdzwjlV4y6uIVMGJAA77v+mLRdNzRSHrZmsJzX6YInbfVPBjRd4DoBjcE+
iYwgau/Sz0R6NU4qBr4dlPJspO99FTD9YbY/1N9prmfMbYUft0KbVNwHh2g/5syZ
GIkUtkoDKCdALu//q9X/Xpcb/O5dUujv0J/3OgVM5ZsF2x9Ht2xKevsnr8B6bpqP
E6yorv2hp3SZfdiviX5cf42LNzkm6WHiPhlzl9xUKHFkXN/wqyhgMYOuh7uj61Y/
jg5Y6zl0WX4sbNzh0wKJbfv1rVUEecpx5RX8EE9RMkUrPmSNp8nWscE7W+2T+I5v
3fqA9anW0rha1MkGw6v8G2EnMI/n2V26CL04E6rD1v6nB2fS5YyJv/CGFKs5jsX6
YYIBqAon88EFa+6qk1uBrQMqLOlRZ38uwSoL/TZDjrwDzo2hFAE8lkMu/JsJDuLd
C8uswynC3c3OxATDr8FSL2h0fBeiZHw6E080MO04iDtqPAdYfcf+BhWJsF1SkfNu
wgZdwuxLWeErYu3X3Jn6ok3UVPYdUdbGxQsC4wd6YAjO0fSOTgBoE87e46dvnYyc
47hh8BYWoEXQUxJJ1CvXgEA2tmiALccSw5ojj0zdAzzHETdNE1nuAx67TXYFeKXq
YsBFl5qkA3Jl5/qFOQN9sfJCTqkjTgYm4pYT5Pj1gvpeqUe1fZtcLUIKWBbbnrrw
cxxn4pQ157kZr468MAstOp3B9a23A72VVYjVfCK+r6neVRYrxGaecAv9NYS1ml02
M//WY7DgzdNscBVMCpMnmQpcEEmCkAP+zEu+5qqwiMToMb4NZGjsh6gW5J842gnZ
iYKmwaE0cdXjvmPROKLgPyL6dnMQrq2PJuMmaDyIL+XcXOyYqLE24Iz55lNCwEnz
rbSDc79LQWyaMnSx9tYXvzG4/OwIUaqasNf8kdCSqL2/EuS81cyI3zDI1JCT91PY
zoquxERLpoxHqty9OJ1F3r24z9koU7+x8ewfXivWMWhpPLRz3YerAkv7CwanTQKy
Y2PqvTEliN6YQZ4yi3LcIKNruwbAh0xeC8FK7R6Szm8bmB7jaGxI/LaeAYOk7FRs
6vR3YDLjUO/NcyMeodwx/GrJRPb3F8cSmrne80EOMtpeWeKAQXyKoEt2bxFWQ8k+
iPdZySAmFb6D9CAhSHeR1F5obem4M5hnred38ldaY1xvaAnxGPa9aV6OxheURFpj
ktVz6DILbeSvfRf1yskirnekyV1F5e7uhyfAMFqeB+iIEns2QRsks9ARyKj9OPrf
XZYXmhwO/QgG6sUZ91KLSb6ZqWwd1aFzAgOUfsFfzf4B/iofPb5zuV02uPPDK7/D
hbPbCwOiph5Kr5YhpnEYzJCtviRx9RiUADRfFMpv1L97eCHL0YuS/oQcFSRQtsaC
EVeKUAzY3YZ/OL0eofe+hbUe+QWovp7Is0wDp/u15eSbLztwodSkGHdggkpO0Udw
y5EH3U3fYNceq3HTaKc/kRMLIHheLBuA2icYilzaY4SlAMkF6VsPF1JV7YA/pz1Q
jkW4gFxRoruiCBuEmoGRuSGR8ldmHRpWZ3xIUq6HzrGfBGzPJVrMH42NX1YSa009
4pS9oa4H27yRf1oOkLcbPSZVEmP9tP7Xa46KEXKCbnfUFvsEDaNCkKNXbxvTEI4p
EQnmv+vXrU3wNng4YzbATTSLdMu1QSHjT1hf/7hRjbLdc4Mxmb8+xOhqEdgTzK8g
/ygVbSNXIpUSIMgqYIRZfN2Yqf4irFw5AtgJ9fe5YxPFGvxRI+eQ/Rzb9GjK5sGk
dLdypYQBsZ9P1P9hfzEyR2ia6Uua+CtHWQDYBlYekgvIkgwxtatKU/3+HD3WM41A
MEyto9U4yidyPxrvqjw40N7RwUVnqjFFUvmeOuOoxfTVoAqlC8htWXnEvXqkjIaW
TQL7d086BUQ51TTArqX4x37GwXd/IhkncDXPjXbgv3TURVnmXM6oWuOks09URW6V
7G5Pbv7vWCUVAKV5bfkBC6HmIjVXYHxgMmpqr5XbDzdCVFgOzgzCFgMUeeQOB8nF
NREgpOtKxcV0/x2dQY9aqSLREoduQxR3/a4ti4pe0oxNJRSnAKOOdrmDvjvytIgo
cImgof6r47pdibo1DWb0stA5UbL1GP3Ez4eC0obHYI8K58/aLCvlDxtJjbMfcV7K
oRcJ9nUOoqbB9Fg/BwDGhfYr7qVmAnz9yvbc7t6BBhxKja/+kRECwLNYm6TGbBjP
zmL+h+jFzK7vJRYRkiK2tIm43+UIzIOLOI+adKbLaa0iUyGglUG8TvqcHunRT+Fm
ysro1Ly9aZhIHCbg7lLKMBVorevheYLmYNirx5tEyt938MBko5/jyFf62aJlBvbl
edcLSsEOUzA5SLs+cd56gnOi07gHL01Ke1Il4yCb5uKZzdXvK6BafhGMOCaBsdcl
a125oJp7cr+PKCqVq4kvWyb6lBVp7dpMsF9Hqega+XOci2Cufl6T5ISx7pW2Zaop
gqxFwf3nCyG0uQ079wV8SE2+c5C4baMZMQTq4TLGobZiE35Uov7Y6l68uP2AMioL
SAdvH83Hkkdo0xXQXq2oYrqTDAXPvzRFYH53aFokWize1XHdWecZjvHj8B6rS8NV
2d9afZ1Rc3TfGD2ncGRZfM9EXdW9Bh2E/3GD0QMDMFmjYbPiLL+6VRo0xcKuv7/E
Ne731p73UE/vejoDcTZfCeHpWRMfl6XZ3KSNNfCuUW0EDZnhSQPmaAEXY2eV9LBS
ebOqe0M5p75xSaGz36oSO/hV2cKdBbnm4e4BlAv9MjM/igd0i3yUGOIGNq9sgdgh
F1BaEJ77kcGSpN3chrm4X/mj5KiMlXIsNB3tbeoNxO4IeRl4jdHjfd8lHfTKdu+E
q0DZsOZ1TvWQkw5iC5sSZGyxCIrF5FnLm57q7zqVNH+b0rI9Grr6rNQBU36N6pRM
VJi1RR+GyAEZPoSo6iEymqB/Y3i6MyqMrVVPfs0iVbM3j1Rdl1yor/f7ldQ6RhvC
iiEkzxo7HMP9ZkRgAgGB56BpcRJhslrZHYguPQAQ5rh7YCL9CSquPDFXuk8y11K3
LdW/fiv/phu1WKR6PbAATBvA40cVRVoI+kEHqBWt/oMDVxJbjH3T1U5oRAMzbEfs
vM/HyJkb8sg99cG10GWpaz6Yx5fk32HkrIL6GjRsYC80RxGvrOUtgqIDcB1X7ysP
wyJm50ptdtz2pVnO9nZABnE5mQ/6ttTsWKoMMm5Yxwq+XmFyRvRVUL2W/lKQBatl
+GBMNFaOcIdbYnCAjfeTjMg9YPj/n32E5la+uAhkkzLglEt26XbxaXo/y24Fpf8G
uaXz8nIDdr8vb/kQHTixQDaUdOG2gbytR8uMLff45oLu7tusi+mt/Im3tdgoTPfD
/9L2zb+GxdEfkMlx3ni7yHdhwT1ROUU9PSBQJSiMVMQAL0lvihuhlJ4dxBqnuKgO
j2N5jF9mTIuDl5K+TP9R7yPIkqOyVGDD+kWxE1qd/qKDivgtgke28vMeyDUyMYkU
OVBXKG5256CiSZdbv8k/ImuOWezlRg1qqJG41dVIhs6PXnGoEKgD77KxsRFaKlwx
qw8cK6xroYjMJHqP/7PMsQHcMvF+6QPJEXmMLAiNtWFi+jpCY/oqC7nLD7EshYit
Z2huRvpP5LP27pVaDMtVBdhrn6hUAKvElR0Npe1xv/mdN5i9cUTAbnseRShXjDkk
9ibhD5DyFtuiXeouBTClBa1PaH70vqTsq3lNqgSrv71jbSwV4wHBhhyTo/s7CGXS
RNSOntQfS8uLLlqIWX6/Sy/j7e/JQ3WbTfBOi8Bq5RoJHX7wx5bPrS3zy9N73jDy
XYFgeE+v/MteHlK7FI81xGbTZaCqEeUDZ1kaGkOOOtrSlvyCjdrWeI13yxk+Ybmx
E8usd0PZsXz6uU3UFrwHb0Do1dRWSldDsvSrqThhFpyrrp7tV851m+ad0rzcKZU5
siVbIf4E7oihUHvy6BPLoQabaXbJeBBCdhGsSVggmq5Qvoj5h/Vy9npQz5RsftLS
ssHzznjwC0Lu4EevSSmJ1xo+GXl3ToO9qkAraBC4Zq496oKcCfzfvGIb/ftXz+f1
mIkWq57HhqN07eyXa56+a07FMzEBZJ2T7bi46lcRJ+LCx4NgBO0JREzSMcVB313i
Zys1cJCum0hDc25rE5c0N+GBEORWCYZjPT3Key+n9e8rIt4b+yG5nE3cENg8GRA5
fcMiuJgltj1ZNATnpYTnuNytwISh+fHvGRU57rxzVS2YdMdYyoCXJb7tL0f4d9M+
dv6wnCiORhCnnJNexC7NXWFlN9+mkwevT+5OQlP3f35gSFlzPivErUzHguc1K/Hr
4/ApSQlMmDeaXkhyKg+rRCTPOOAjCCQW4iobryem0zbZJwfzJNPoq+nZEEe9O7+z
YcJzl4ZkvSnwhfpuWQiKCM8o9DToYufHBb0CjWTi6gJoTbLpjjznth/GthJqkLZp
pi3/igvBYq9bA8wf9M0RPw8xBHW3dj177LmMS7Ra3AHfpogQLMfFnn3QmS4fKIf+
5T2gEt1fZKfzU0XCbsgnQDsmxLNxAwNCfiFHcYcbnUfJfd5rnWAC/gUUSdNZslmA
4KXtljpXr/M2lRGtUkT5fJUdY3Ho8EOhastsSdxmdH+jfvLf9O2ByLAioEmoXTdO
C2A4DJ36T41MnGUMyuTYqjJgkNZkrD1jn4luIsm/lxRHq2Esfuc0L7k8jwMIw5LD
5i5xirV6M7i+FKzkxmYKNXz+8eyPp2Z1y/x7Iea6feL1yOB9vf24hkqvJ/UUXwBk
j+PvRgIvRevRImi5hEuXC5H6zF+6fEqU+4gX3zABhwJred+5dPJaAs3zRVm/h0EX
yLcrNXraVhLVv054TBtST+diehD8HRl3ZRIgjmCoKKIVAqW3YVygRe3yNtEuhSGJ
GkKQA/evFYNuto54Ttgg6CAkAIlG9dUDVIBcJ5EpjPsXZXYHolXq4GYgg79aJmcK
EHyebZ4xRX01P9Jt1cga8kjsvENudJFS4fH4IsghNQ4l81bxS8zdYqcNIgTXcVkQ
7F1G5DNThhfVuwfYxZPGTpQpNP35XIYIg24kRVgaU1dF5oanLjwZ2tM1YRpGj2JK
Ameb26YkbGwPa7UuWWQJX8fhoSUaXXJ3Abu1Ye1QJeL0Fck2xysGwnkDsqb893Dv
AxjTj3NQXQRMU/nLpYRFp16gk6tJrJR9sOM8w/PJl1tskbKEqsEfHcZp5lqW2KVH
Lgx9YgPsV+kSokaYNu1zT4yS4kzzNw+vXfPt7FDuRrbeIZysOOFfXSbvFkg608uF
X3EOqna084td+aWHcBhEpfasJ+nc3bcm7Mx7HLjWtWDBRdLx8+ionotsBMakb8hQ
/FoHTm/LGUEpErpDPwtue4hNo9V16EL1AuQQ/7pBRZyda7E/oqv33BD67oWjYfsd
0maNHgKQsJP0Tc9MxNd+yierMC8Nlful7Tt5Sewe73jFRf2CxrVPkhMWyVNtoFln
TYjPFeO3eUreJJ5HZ4jWtFfs0sUDFw0VrykY72nc+cfuwWk33oIAAud3MuLCasRi
Rgp/N0RkBVCk3RUkncZCRUsP1tme0IsTaqliiorMq9y1KBjcmd21jmsAWsCk7zBA
VPNa6T91IrRVwSUkAxpHGr4VpL53I2d5Rcta4SMsfTRc6rt9bCrn02Ziwy2aIEaC
mT/i4nP8ysSiw5PL8I96QT/yyTnT+u56SfsUUfIcwPcIIeK4u6pPALcZs+P5AVPG
EUpurb059BIYtdVlusyQkdFZWSPJlLw1KnCk63YjFmlQmn17YDRVqFl3MdMKO+wu
Khx6IMXMl4NZ1OUg2ai2EwYz6JjL3wveGPKU3usYDR/uhb7gze22BXG38xSziHBK
D/AuDhJ4Z7c1IVgcTtarHChBwUy3pWb2AFKbBFi8Zz46jSfuHULDax9KMyOQMvV0
Shbomq1V1K/BonNc5MS+qrJYjvWd1PFiI9DLIsaPw8l3VaX2H/JbJdbj7u0uIvSX
Hh7Oba5VPBlIcXCZAUjlRH81xGpfAOeyLZtHhkmxI22tU3EBLaQ3MttFDYRt8G1K
wfG1T7VaU76D/+/e7dwl4vY1KisyXievgHieofQr3dCtrzzQZANbHakzAaEd1E79
DpSLJnYH24yh2Ts1Db9ostV6aMDCgkM9K2YOY5j7lLNliueaogeeFRHPlBf1xJBx
PT8j19mmyxeWqe2NQlut0B53cbDy9714+0Mkn8q17nqGnMC8eeWvErtZuru5dmCQ
QDDfqvt0hfBXwbIgudIpLRk/abXMoOWNXlT4cF1RuVQl1rysAovFqK7TOBgnXUGl
3nGCTXUtADhW9AyENcRa+uusdIttuKPWX6A5P4UPRr2yiOVAK3MpuV8zV2OQ2xg2
Kt2aPvYuVP5hlFt3KmXnDHfrd79WR5Ra9PirVKWZytrLzbFkc5ChQHhHDxc815GG
tDOs2A2krT0kbPjFtEMclNQl5pXgfmEDhXlSu4NPvhftethxd92g98e+CGl0FQTR
5DNARLLYE7gNCgmGXYtGCXYVyhW+e1RZNoxmMz6T4/Du0zzfP/LdSYtXH6Bh3t0N
kIV59ClLjbu9pFGpFBrgQXoOY/weiIvWr/fxlYxUUpQyi5JKaMcMYIDrO9XE3GJF
oAqgyYbPujnET0T4Q0mRkcsAgECDjEo3I4X48obZdIOshZIx7ejpoKTStv0DEKeN
sefGwfAfsFfxlixYSgzznt3Em6LUnLmNHUYWVb78rM2vMK2+4oUkod5YqdaIbbfn
xh45xCQ8tTpBhkadH7/VmaqDzelaztTLcGUTSWkAQ09W5Yve8ffU3hHm2JL/XDMW
MbLAFdCcWTNHxvcZZpVqLh1mY4Bec2nyV+VqZp1WRPSJTDuvCTJ4t9N5XJwKlcz6
mbrualW2FcxnP3Q6pzuTs5+fmj4MhWb8pJAJlJbg2RTvF1MH3EY3p+NK+0Ed1xq+
OVaARha7WZ8gcq5fzfdfwAixaIQnfXAtFOCu5t0t0cDhzTJ/c1R0+URkNxbiDKVr
INBEd/Y0rjoolX3qN2Mxu0P4yk4dbdQem2LYFqeMWYLTtLh1gjreBiqqWFuGLAKr
bT/2PBH5FQjNKs+jnO/5mnA82WyEfyqcsWPstigTsQl6a6XnUIEL49F/YcFHSjOP
Rd1/15F4zXyOQuBfjzGFKynKU1DJX8/XMy73AprASVtvzNWVfY3GxWf34wUd8JW5
MOSwstv3XY1qA3dI6gdeDkWIvhjbrxPw56NvXO8WleVejXHyl7tqZY+LrDgj37qb
wkEup5XrKAqhto0A4sWTRaFpRAFifYbM47SWGdNS5OYl1DpFwNk3pRzXqzTWxGuD
bdcm6IV7EXkuEcl5fhXGZSUIZ4A7jHkQaeROHfQL7SkcFAYo/vBKr0bZwf4piBGJ
e3y3+GsVkzwiMzhXZS/e6zDk+EA9Vo3oiVJEQUV9/X2uD6h1w9pqrUzJqQlynT04
m8wIlCDZYVSB6MjNIcPv+TvqqxGvdEbIFFCyd4ZLlVoggAGLouMt039q3ntZ+O8m
qgMVz4epsV9Ay6OYyrU6VWOVnpmmX96Y6BA/arSe77+BO7JejAUmanSezVtuVHfO
dAo6GkD5TuLxgUaFqpnQuUvL42qMsDkHbzjll10gzap9Bm7cCEjR6S83YaT8o/dq
Mlbw8gBnJyVkcx+jBiSesw6ZongdXhY08avvOe6bOK5H2K87GJSux+YSyYqK1KPJ
y1ACJ4D9p/mLsaCo/KJ/RWVvhAKqAwV7kM098iMAXgnezvv379LmEvtfUINyWpju
gQwngHbBohn7A7rIfbEf7wl8MoKCN7qFyxHTDI8unXG+jDxKN0DOG/oK6ky+2fQ+
4hk12uxVmU9+Yr5bHd8Qrc4sE2ZHPRUSisHPToJJ/Ln4954j+yJ9vqQIdKmIkXWa
YkhNRYDR8gmcIop8GI/oQ4Xltr4urnOsivV/DOUOr0ZKnzM8rocppQ2tO4ZskTDM
I/Po2Rvc/DtGwRjBKUhwJCz1/8Wz1yaI0ZeX/7boXOnD8IgXpteQEVH0sgA2nhsz
p5Xsl4oR9pyLYnWgKFogRJKrgqsuw2WKJ2nKl1UgzraFFqemyh6J6PQzAYQgkUKv
FlHbOkApOxs5REhMczcjsHciiQxH/lDUtlCZGiwZfLMLOvAQ+xlQdAUYQx8/Esn7
iMckM2Tsyvy7stzrAYU8JNymvWZB6s0LW16MfxrXOxjnNgoiX/aODK9MEUaiv3ow
/d8SzSG37IezfAZURNGA+wNI6BYKXI/9k4GkYTvobwr7lE8dAJoD1DkK1IoIrFMP
Z/pXlA3SL2nwaKHQLaFUVSF/LlFQbkjgX9nXzaCADcpS9lKEIbhfv8z3FaRyRQR2
sPVkRC/r5cDtGfesJcIAuk60nRRyvy3sGYXlh7JWMcyCrQnWLLAataZaKIrXExN9
7BiT6VsYeRjCz8zAUg+vtk1qpycMDlNfz5ioec6u99d3tAHA7wr2TxWKZJTDvLtg
uOWuw9+2s4c21ttWPprmHLh1gLUXqBgaJ4SjbgCThVzVqcaqBtt0iZcmJPmv+nTW
Rmk9voz0SCAUGIWFfNO8Y5dvNtXwq4klXDuZgxvh9XS7e8S7ZqrUvXljNZLAjc0v
JH3uepMPTOmJh0fLqnDaEHUg/Jyla1+F/PImJvOqjAkRITX0n+KCs1v+5Je1J64z
b30ast12HilT4P8NsrA2R9QlWPXwNNMgUebLsyt3oO/vjw/T+PF2QphTQ+HTv1Kz
lKS7TOfQ/0/b5LhTbkbiCmFswMR2Fbut8Jj1R9Kyi5CqjWsWtyHASXn5a0EAwCq/
9Q/KdzAJb+Con8dlPa9eG4gpp/orzt488yE/AKlf7/tumGi+fcUmPasDvBBvvrpC
I6nJKPETSK4nMwBO/H12J1ynqhTTYsyUvHgLurYvrMIPxr4xVh0h5ALK/r1Ytg4Q
+NZL7QgvB4j1tkKZSgO7XYP6878JfLAOz52XnAjFz5vsUkS0RA4nvJ7OHaspM2Yc
tt/8B9P0INAFJ6svT95ArLFyWbA2/y/ne2N1aF45Ku6YGUB11cknJkU3mHZkuloj
Cogb97WszFyf3PA5ztBM9+qmEvArYvzA/SrmegcN6/fzgzLorRLi5ipsNF0SeNLc
HDaFeBidW0xx/b2F26dAf5NMVaVDcsw9EDhGb3Znk+uY9xN1+l5wNecaxV1sd0XP
yxzgbwRIxiPjPK2gA52DcyRMWRTNAIZGVpr4PG1sjIOyp/zgp00Ag9+a9V64LbXz
B9KILIVi3Cr3jfNdUKeYCdR02hOFjrHujtCltvSEKmakDbQ327nyhWBvCa51VYhw
Jnv1pd66iljSJGQowZumiXuuDecVR4vRASQxWcs7UhPjmZwKzBah+MoqV8j0T6Au
KIo4oJylfIxWug69t3N3vd7qbwuLRaxTGkUyP6XmLiNM92cELjwAyXxZ51cGYBsP
pwKG2pk12cUHcQylTSWzEk44SeocYw6w4A+p+bP8LfT7NjrESf+goTFl3pW/ldPI
dWdTOxSueyO3iXCjhz8Kz917MQrtMl4q4BiHAVTwR1vSFFd93vrv5cC8v8fV1OKF
Q2ITUs2YH2RhgEHZ91aixusnOIAh/6D3dMeh/8LehwN36RwymCB2sRB84wkono3O
bniI1oWjTQGSrKgyAYwkzfr3I1XvbpjY52t0VT5m5bSJqU2hWd5DrH+kVQF5ky/x
dySL5VBD+h9EFY0ra51jpBZD5iDUx9GlCS67s3DvcAWI/f36fyRnabfLyJ94A9tQ
3SHTZms0mmCl046lRCju1Gwz4FkFH+uHy61fWAzFOSn/EaO/O92/e4g1/vt+riFB
ZwiNUvQfWb0ee2Np87yg9iubRBdpYPyB2ioMif6VK9voLDsrwtH2BWySXIzMlkMY
GAMZTeujnYoKJPoKhO/eFMwdC6yqX3y46YORMHHmBB6wMbqKJAVlWB+332ClnKub
rM5a8f2ZA2uIYMLp/7CaHghF0CUSKoa70RfVsLQ4EZhPYyiMburec//wuC0EsCLE
eksdGiF+HmGxSA7+EtgYLpx3o1GhXLB4rY9tjYJSVhTO8dQDC30xBHzUw58l9EtG
GGYgoQcpdsNKr+xQl+VMOzedIHHP1TJjFI9lkdE+4jGNwjywVxIFhXgGD0eeerxq
/xrmnNfXTSslyhidkKar5SWr5g8A4ut4eeqyajPOzAv6wtMlsBrBEUXL8vwCFXRK
iUKzQmCldU9tk7fLkHM4gM8Q+JjmkZ0vewtl3wjgrqmurAnOQA8SbhetumHA78bu
mWcfmyEJbCR8a2UlKtsBTAEv4W58+Jxev6rjDVUpLVr9fLep7FcmWJ2EpiJYgLxo
zDQ9I1DzvtxiWu9Poli4n4QsMQmgx/6uVl0NbCUN7Yx76nQjPTsKJEBuw8sWCIQQ
nfT+FXrdzEobyHHoVWqnPgQyyiudGKZsGAMzNZHBSmGEhKc63HWug7ZNeLINq1zj
4VZ8MEkQnh+UooGVVLM/mYcZvzAWNHpAJpyL2zJUO1gShhnxvpQlGH/nk4vkcZf9
a1lN1hNgqAWuSRPNWqZAAHwNZvI0hDtKd20Ebx9CWECbEyvy4aSgx7Ht6J0TtiFD
JWnNTqZN7vbRAa+7xGUriIsS9QflyOofETBN+0LC/2KN9zxHMcLaShTJpZLnreKW
Dk5p3/nVlepTED6ksO+VkZMUlgyYgzee0apSYxeZYd7kwBo/+HBqlq3+ua2oTAme
KxPAA2A8N37saSoNALqmnQiSELMveqfxaUxGKwE00TtLMMuAHoet2bB0+YtzoZeV
a1+8S5LWjpU3qwY5bUnzn5TemE0L/US3SsdZqgTfQ8RX5aka9Cdk9y7TSndRPnmq
aGtHroGePFgL1QxGg1iMgolO8pQOh+7ISsToIbIwx2awJb9mljSfoMqWkRfdW2D1
UcND4AscfysW8/SzybcQxQ8kfcE/oZ3z7bxdpMXj0AnSft0WmPXK6BvPAD32IQLo
m+e95kDrPpLHM+vUqnnTo8e6v61Ga4S7gV2kf5nsn2kXZrhTR2vyOjFtiwJPFfXU
fPM0B3n/CaDeo0Nee2arDdxlYwCCFiK8fjrrZ3Yy6v7yWzLj4UCFmJeVKVMjzV0k
usmegECqxczamozWQXHoy2pEFb5l4oYBb8f6h3ozC4/VPGZrnXXKwH5m9m/mI1VA
SGKT52fwLzE/Fz3YKGhUBKo4b6jKSAj93tIm9drUMptYoIzOyijSIb9qoThPKGwX
/Q7PlAyn9OW+ds3JgpDA5gmwp0R4sk187TbrQ1dd0HC8lFGKKPM9VQsDwV4NRbrF
NkllYhq8sMuKU//GBQeOGOcToXg+i3zbEJje8vUVAMUAaCwBpEpmSXWUzd775ARJ
T+AOJzpEyTaA6ThMHjyCwYGRxXiw9y8a9GIu0J4uE1CpUwQpFhEeQveHzk9lKJ4C
To/HFprfKhmOBgiiF9xWY0hxXH/JRznh2k0Wn7vTBj2vNZ1ghe9k4Htq0c2Qfw1s
Bn1vwzmXSngc6RNbZBGaSvtShZfosU4+kvf4L8031I8P3LeRJFkUjF7IYBOz0ZUU
CAwCFl8YVgUjpKhR8YKH+R8vhu2alFZj21e5e4bJqnx9y2w8yGDQ2AgxBOwdYGWm
kAbQ10dxr399qoptUKd31/bW63nUrJyzj0cgPByEpz3Q0fsY0wW5LfCAQgLQ4DNm
YxI9LNj9eGHQwSM6JWYQIpH6AS4zz/kWSt5L4mNfJ0dBK8DMzP5P9+NV2/XNBXm1
2IqVnRwi6PyDXpvhTL7ifmtZZDu5/Wj3Ws0ufXncVY5zGRCLf+qpwyLeNIK3AptQ
f/GpPB9taQ0Pb2J9m7rNBEoK/M5LFUcurVXSZxRsdlZ3yhW80lb8JbO8KzCWONNe
g/0ccnsDYLmLDmCzvFs2sfwsK2I6f7cpoxX1uXTkyyHVVfrstq6Jcq6InrOnaFRC
jbZqkNVHtMv9+D4TqGAUIThgmq0tNH43faAOaK4w7Nho7nKYDnr5pkk+KF0+b/Xs
IHrbp0DM4tQPdxNDzABoXuRTiE3WWlHZLP1+SalaQ2BQuv1ZEgv4NdMgrIRApQXj
jvnqUpl+60JiSyDzthpxKtTaHA9AsyMNJUOVi1+9ezLC7K5SZdT2iGSN54lnjhId
R6QJvCbhlhE+6o7qeXsFbynBxpC3q6b3R/UT9kNH6GBcMqamvyGlONoWlovOyWLv
Y38HB0n8pONRWNmnK6QbbwvWYmnkBKhBZXRW78tiEs+hIH1pURYiYn2CQmuAs1ot
tmvDp+f0fZmLhMN8VoeVFB3lQ6343wgjZYP2zESpHMcxKUOBJfEjOwrZFSr3EnDR
s78zPif0+M0mVsonHCKqkfhHsycT3EBnSXLKg5JNLupKIW5S1N9qckjIvHssz05V
38zOG3oOORkatADAji0k+595W9MODrX7mgTNpeckQ0pKHoNRBl5be9GXV66pSZFa
TeG5AimlehPXdb4so5eiea9oEa/M219+8sBP1ieeO+jEn/4l4tkeOre1Sm6kdEjS
triLF/iMarQbwpoaMrICYF3QMogJsbBHBrcS3ldjvaR9CPIiGr1e9vwiXTVg3+ls
SOeudUvcNQdj0y42rMJBcQazeRfZBlOygkBUTlhpS9XpB+aUgaz+1GTcMhhXJ5TV
fMdlsGwHsSXDlbEcom2/3WYSyx0+jor8/J4Lr46IV9YAK1yWRisP7Tz0U8KBCAEm
9gJjY2JMBfvgvSARnWpu4In/BFZd/YRvz7AS5XV8dugP9hfHvyt4hjFgQlVxNqLG
m+AdgPlGp7XQ+7Zj9+Slcl8zdgq4751Uia0oswsQ/RKuArHZqlH6bxAfpFGYiKBR
esST7SEWo5hhlze0UhPG9b7t6OH25hSAe6Njg070vCbbo9UJ92kUb1Sf8duKYTrW
Jw19DBJq46xxb50x3JGw41QzBjB3l/jq/PDBwUKmGtq8QfUPp2HpUmUV8a2fcKDj
uMwIumDF+PpOUk/Dl1M5F6FYvaDmViH/aPr7cGQkDcus+XXuuVNzFpfaXdhbaN4y
PJSD6VdWizBIiWZxBKMFY2wNDXMPzf0+S/sRrv1smbWZy6NZw1H4CxJs14oKph6q
P0uQt68gVFyts7EMRh5rjv1o+kblGeslyMlEOdCHRJrj9swXeTQAPdWGpAJFNTeJ
JckQRJv1nWC6gsxZcFT7Rsj6RbBHzXxX+TaQsZXaN+Fq4pj/fTY7Bxc6GcyP7SGo
JQXqcBZihkxSdGhupWYOd6SQkCzDL8j6psqVGh+shDGTutk6brv0k5tC+yPIeckO
vYdHibzQ6u3l+AntMDcaQ9TR6VRzD6R2SxZkMsa9+TVh55rB2tbVk+BjKt5oT5iD
4u2kyM/5XU4InqsU/innrnlwnWwRshPI7BsTG2cWwrkX5hnYg5dJPkccAS69HnOC
FUvFbjrnLHtFTl2pAsDrhlrHyjx8DAsSJ+4GYl4a4lNhrGF9vTB7AeCNdNf3dzxs
CkpMw2hkYK9syUDII2KSnoh0YgZn1wmhwWqeMU1pEuHHeG2u88xoaEuQ4ctseYiW
H32sXqPm+5ow/VIbGZdxP92/V1eMVjvWbsOdjPxxmggn39bLgEYz6YhbO27wI9Jd
rB7i/lIsklP9BXZP2oeifUy+3+KaObd5qH8zbGqMCoBveZuZdYZbNTMv0URRJmUK
DEfKIo3nRXrDV9XuIt6ne46DBe+xlK53l8+iLJPOmmFuPlXVwTQQSihp4x704BIs
POCtC46XFsKnDFNhbYquHzZU5SsdbB5fa450fyJKyQN+hvfFg3IirWwwYMcoOEI7
7grSryjP2iw6WfiM7JF52JnQjo+mqg7xFihTXZdAfkWhyNlCnotQ2UavXHFVEUOH
rN4XLKDOSQObbizyYt58wyyMj1J4TMqRNQis4HgzxuqJbQB4r83kQhhh6TIuApT9
WrdJEpS41wtCEagbEpnmiODEQ1mAQLHlXKnA9aV7T30woa1rFlTwqObzYvLT6DFP
BQ19vjJlRi5tMAxLJqyW68Hb/dGY29duYKEjRDy4t20632ibSMzn2hsvHVfuQiIa
oyLNbbUqYERemdTdWMrvve6Styros6kVdY2fQmq0DJ3Z4H3Kci8jYnSILcduPJ3z
VyH6/CMWhwl/teirbbPoL0c1TzxqaRzQGzNKYXkYXTduRhRu3vSqpknMTN2WjUSp
kG28bpyuBaNtd5GPQ4aH4QACFSoYBA3xCNeFlqYvVE1c5nszgOf680SIiLaB92k5
l6OeMHEyo+2RcMUHhS1Cbjeni/tdh1za97YFWaAONsauUPIHKw1fg1AAkR8xtqNi
NaWdIz2q6bdkdDeUa7SLLqBy6N2lAWHVJ+lXFoN02OTtATn64pHgUXjTED5u4B2I
qx0WXxKU1wyZ3BwOIZ2cMGumDrkcZZV7NL7LSgwOZ3QHD2y1MJDVnt04w4E2OtH/
a7c53tV8sMKw+7bKJGIBBiJWUdrWljIOdktCjAkEaaQiKF4TCaIHOxx839XdKaRW
PHJyNitsj+GVGUW28kyh3H/eP1OBghEKmbTTVl9vjYzOBET4NdXELDOXhPaqel2O
oQNGjFyWiIro48+N8pF8fRgEDyXVBILjb4JeoJCK5X3ELfkSRrOWeV24FAy87Pj4
5bigXl8JXWHDYAUOFOmoWBrDtsXBgrcnkEv5Jmdjj/DUCytrPZdrc5qUpBtskpyK
6+yFvFmc8lN1zEOcyO4Y94ij1UVekhYKIS+NZ6F/RQlnD6koDXntpfdj8GHAGSzO
DMbpuK3xAkxv5DdoXn23pcrw4s197IA7x9+lFav2Ds91LWVJFwVJfGRZAx4RB890
XWLfdLMdfVZg7nPV2OnJDoiHZPnbvfk7kxGa+m3Rdmh42ETYOB9M9uFh3sEJ9NYQ
VZsaLfVNc7poS6E/iyUanq5cDnQBI0ATB2mzvM3AP3FGfWrQDpBNhiuAlIJZlyrt
fJQ45X3qCs8ADDLDBw4EEVpUeWbBYYICCd1duFmnswvj+1h0+MULy5pcdOGUrtMT
hcxibO6KpoO5l8L/hAID57SWYwmX4AAJXeK3CXomDmKtGdGqUalf/0I7wi/wYwzZ
GXZxx88r9sEBUrrKv7jfS6++rvjWfJvbjBZGVH5qoq5gn06Qdp3sDolXbw7biIA1
IEukcZAmfAAaMV+j3C4KfODXDCxjqGVeuHld/5iMAr8sv6E6Yn2ci/9zV9CxfScX
pzfK2x0YFD4VAbIUXFMPwDfSr6xsk2Dlk6fa4d9GE8NxoUYTRih2QIoHuRbgm/Pn
N10AT/o5Dkz7pGvOZGOMYZy4y9hPk6feukXs+PFOi89ZvEEYWEccHDyLwZMwk107
llmWrdLL8AbI67iGCrjUUciOyvx/0ZCu7WO/jZAUcdw0uceojpBwH3CWHuM4gmTH
eFW+vRQX0pWDFs736mitZYt6r4iP1T9ga4N3vg23C75fYnDid9hrHBfpRw9KaZN5
T11wW3kvTa2B/GMEDdS1KlTgYA9KzbyL1kCyKyr9KKu4g/wsByB9eNAplMYifxcp
gv6cLCfvV6jmBkkQ2160D1cQxC/rSzeMMvjeuGdSRY6vb1UAQpPQTalF7TS57TIA
q0dR2G2d55xy//W4DjSXGc+07vUvzZiw/+S1MYoYj//ln7J+OoAvwY9YS2aKuixk
jr8UPL0M8uXXHCWDOrwPVpl1k5edzi0Dm5YwT9emY/w6ghZ6L0WmeHJkgAx2P3Hx
dL01nOp3UhS7u/T41opAV7wiTgB01L52Lj9xEcGgcrF97Fpu4poMSKcyE0/yNloE
Ux1FQtjO6LpE6RRa42/sxlrv/aDUhiSFKRV20mnP0+dKNd2AivrC5vpL8Jb27C7O
ZHF4OKo+ZcVV7g9BFiuxo/51X6aEg0Cb+Aq0VPX97Qu5cx2M0Kr6yo4bhODe+ZSg
BazJ5Tij/IbIexMBKa6XwMBFI7Dg2slpOch8t/vDOsOWqEJfHxR+jUIbNVGdsGDs
LMLN402SwWJMVKfiIgThV7xX9JB0Ab96gXxuU3Mzn+f1oumn5rg92lXJUZnP34V3
l96zABeDZOfVdx++H5fQTNA5wDpFWTRjk0nBmJKqXRPjd6s7z29pcPGLMKmHclcP
s49gABBo0PwiG3LPL7A2OS+tD2wkCtIv6SxTz78gSYbTPROmSq1nPMWcwh1win1k
iEq+m6D3W/PyonyviC8bkN6TiQ4CMouQbbjI3+WjMteGJCww+m+5ZO8MeYD95rVN
CmS93ihRJqbn6TqlpLnQsTrGUS03bjSrTfKOin9gfoHn+7mD6qYWQcHs1VHhxFoS
Ra/neZqZtGsku/H55EV9hg5QnPpzVHILorSAk8XQQsuThCQXQhibX5bu3rjBofJh
cF3lTJXArVTyucBJQ6OynStFWRp6mSwagvqc5K9HiCZ/QKHLi2vXZo7RRXxWUA4c
2odPSLz3ErbaNLEIUgLQn3SKbDPlNztB19NswkWm0gBWt8sxw3+svWTBzABVIZWo
tcK+qUfFG9YPk8OEb4T6IEsUIcSAvp+03qqBAVekf+jGaWi7kFP65ImU7t5o6zSw
KZ/PNuTUhCB9LimDW/l/gC05Nc4jYyXMMe8W68ZPkotFBHXK+8Vm9UXL8MGuvGyj
QVp5q2uGjUCWPm0urc77DMcx9Y2UaNBqEgJbM/wrZGYlDCj/yEUOOAYnNVwE1luk
edTG3YEBkAkbQ3HweQySwaPdYaPiA6OZ2mkwcqgV7fEZA0ZfygoEYY2ngKHoYduo
wqr8gaDg0NBleLV6A9sIl5qKLLK+YhFNK8G2bZBfAJxj4W6/ZpkRdWh3237VSuZW
U8/0iehdZKMJum/HHF9rw8F3M7Yv7FGdTEIMuY3BwY+BEBN82aayS6zlUw+nSH36
NmSawrnig7aOiSlqm1lQfGbCM50mxX5V4KrFD9IIErbGHDeLZbT3sZIaiTmYEeKT
I1TBegZl3KebCqjH5c3heO08qxjMfNNdMRDxG+T0zobDOe8Jx8C3lTv/Cz0RcaBA
eWXnt3nTz+JpLIMqRIjlgwdXG7Q6Ast5hl7ie7bcM/Yh5I/MH4mssMNyXJDeL4dd
ulEzNAqLhJHFX6DlMQTqBpDY5X7zJxSRkXCgSGlNy7tF9nCKxIjzEBPCjdTkhBZq
xKPjfdErFvVsMXwyxVIYWc8QHFpXqXezC+X+9hsJqixgniwrKy7Y1sIaJ/ASmpQH
lhW3Uy9TWupR/LzH8WX+X0LeCiDXTQiqRk7lr70DsKSXALWaSYl7NB/fe0xfudhE
w1/0SftC0+7Z4rMXHDSCK/4Ty+lE0uD+QxTjG5df5crI75JQUuCyiWab71JLms/9
bxxqldGiipfqhdx8fIHSlBVIV4j0TUDtNBS2VTwLxekaQHTzWoIZDIz1l+Q23tlx
L1Nxc4ZVZUZMJ11gzpHEAQsXb/O7rurUUQtjO9UOOIthwU/AZT23ZzvKqA7ul2y3
jrLQjh+Dk0/8EMbboL/9DXq8eHlRdPmT8TNTp+8IS+8cM595x0yRMPDULXcCzIuz
bITnKhlBVYfPOTwnrv5JtKVGfbjvVoaqaM3mKlKDkgOcrraYKyPb48bIGCdE3WPJ
sZJZOstwRVwU/QADfyXeO5lPY9GDlEKroAzstk1I7xQrdk2IMDMuifMtrpZaSFJ6
tCmO7mP9Jye/6hswJfyOuYtD3Mdf1UXFIDohJdVah/xoskMlynJKo/oYqaPQuv8O
E48jaU1WNKDgArI4N+YIThxYh50cQYzvqCdZsF/BTnOB/l7r8rlouDsfGsp8t09t
Jj71fTTamR+KKlpYTM7BwnYrffGPVuNEaFuKRX7yemmHP8cE+DSv/LVbNu/DdPtE
wUs+4B+rKNErhddZMXLKyrQvlM74dHrefl077WEiHKiMJkhH2iSPTFAW1zTop+rh
/gBYLbZ5zoytg7CThVkNRRpVV/Fw/SToDLSQ0TWpn7BwXHZC1jlcnsrX8hoJatD1
z6wn14mnDPM2YfeMboBwQ7R6iuzU/qVzvyrskCz/yOiMYPKPaClYQ+4qUXPj5EV4
lzjHn7wULVMlzo2cbmxYJa7wYkXx+uhmMPcJFvXYgb27YsNI8kPGqp7sZILAbaB2
YqEznRSYX/lvxD+IydVScQza92+nWvoeKM450L6t8ZVYwj4Oc5d4HWM9hNCW29VK
xAOCo1fuHGPGXm0S68RP3NZwy3kOdkFPPQ4NU3ZdQiazwqatJliHncHbRG++Q1is
ARnlCbtYD1wPNbcB4K4glF6kA7GRZnuSUVXDh9iDC/t2YknMNaK9iWlZmeK7Wz2B
/rQc0JMcxeVdj1m7A3YTiBr2STQpGzIschybi0nBj0W9gUlHx1hhbP5akTvN/8z6
xSA5Oee0YFoGLjrlbvPIzsANIjXZsIS779XWNz8WGVMlN34XvEfCEim0H8Df2S4W
Q836yKUG1TFKmcdWne9sIqFfZPV7dNHDI43xTGjmkHp1987nPmBloJKugxoghQYW
h7pJ6NMLZPtd/UtBNL5/WZRJk4WD3OSjXEJuf+gGLXsikkYBrS/DarMYQqHDYWaQ
2uDVwK7NqBG0VDso7qMTIopiisY+I2q7QhCXXcMOOtP0sx+Uy5u/XY4SDx7BnVqn
iUVzYaCe6VjNlwnM46H9KGRQWpAzqpgi5GS3NabUwQXBzbR50XBtnaWPcXIqF6A/
uCYFO7wh/rc/41kXe/AIzUDSuviTNVFlVhXH1ueQWlgmahZCJ2uCwEknZ7Y9CdtF
7HBOK+AIDSxy/l69noDtJVyrospAH6i/pmlBis8YgZ1Q1x+oK7MHz5kFljw6V484
mkzsh7zif7sY70sBLrmDGktzbm9bw9UCWw+IafxK4Bz2sD8sESnW1nr1+h2gMJpR
D1K8mEKXOWH3TlEdiFDKPE4lHjLixmLOm4nAWD6L3XRpqluW0pOvjPGwO2v3aSym
9bIiblUYnL5SrsL5h+DZOh9zq4dUtCmF/lF1AnAfhvpAi6YcpDGlP5l2jWHOKEJT
3NgIRcNbwIOrSG8roAdhWomTMUdapenrLq8jnjMcTpITo44pnmsuU0cfrx5WU/8w
n+vQZy6wV04iiPeF+v9G7I0P/1wYJ0Vz9fNL70cz4QMtcfnwVnLhklrb80zt0Zn9
k/vxf/YjsdW+aaIyCmvFIuLKIEuv+tl5ouLO3iXxH8z0WmU5lY7fUqOxCub9ww7p
qalvYFPKUH2pamzf7l0y9AlBnGBz7pKmo40EyiOK1pe14fVT0N/llau0CBgvS3rS
QEDo8xwkcc/Q+fNr8mSYjWpraBZS/ZYWbPD1pugnIfq3zvwr3KnpAQFuyxdaAtbz
DmYHLzWvHhmiKUzchIX6LmLwTNacqaFjROlgQs9oKaUpZl/YFrtE2BB6wrXFiHYJ
bfD5Q1VIdPXIC5uTjK7wXe/lexE3yjE2fv6ZZcgZ8H9sCUfg05O4uidj1fpAd/3n
bDA3X2mHZSqMw3PAx89v22KxJDlVNR0GedKxMGlSk2QIfcJqL8sP9LGcqkLOWvbx
4+GIT5+/yrRi62bccFryfBYcGqMaSwNG7tsjf1F1PhHd3dE/AQbh2ELAUA7Si5CP
rTR85i1hm+jD829MhY5FpLtmPshn+qlZhe50D91fG2yXSJJ4c52Q+6Xtds90t1a2
VQjdQNGHf/oR16ucvTQGJf5ZZkj1gENtMAsm2Cdzmi/QVLMeeSFlQtYKzaeUN7/t
mlA4alkgDFxue6mJk1Yn36vM+dvjYK6NuLRL+tbzNWYoRUoQdn3UO3xH2IZA+jyi
0jGyfFTD+AAwhyGKVNKjkNffMSd4hwpwC/uHfPYDmTc9GUr1qNhNiodqmrSikqCW
ECkysDlYt2Pi2U50HqE+tA0A5Zy/WX/e2Mf+fZJwCRgqIJ8jMjI6MOraInlKBOKI
IFDF7P/UDyuCmV6v2zOn4PHnHCUh5bLykINhANYJtvO70YCXSg7IDsRpXOUlmIiR
avfmxpisQXhmvkXdrz5UUFqne4qV7tW2oEJ3I7a53iFVD9wTpl2hkBo/oFZFvbhr
T0uoIAFNHlt/fxJfi+7wLNDYl8GEJM/AC9rmiizNtT9O0fSWgBgr3y5qJNGAVIBM
sXXpsimVVPfDF5XKsAOM+Yny3nc1bA3ZzM+oX8JKXnydGMhEofbkW3cJmMltpF4e
9yPS1lg87eUv28GnZfMC5pqddv6cK4qlWb8gxIkvWhtm0LwZuAL0yTODq9O118hU
cNjtGvgRXkOJGENu18gjXQlUVTCOGbeCOvQTGihUq7Zqn9Z9CR9KEhBUor2od83K
52A4zJEolJGv0T20xZZM6Xdbbkfj5tYM89MhAiUPyPdl1u8EXENHWbR/K25beyir
aiD6xVCOdXz9bZ6aqA8w2cDLaUA35vngJSH6UG2qV/d+MkaTmtK5goviWqHFDNou
Z2GsCP9ZNCAOm4B7bvzlit6EfNAy9cyruKJnLg2/CyBuOAT9jmLQhL2cW+GTILl6
HC43ayFEzwtccIKJrOV/CmeY0HUVlKS5GLQUcJzV++W6iNpDnMFyZjjZdpwkfa41
nYLaxSbN0b454a/yyTDa3nuUWq/JtlJkjLLr27PHU6QP6P13H7vT3UPrMt/Y/kYe
I6tvKa48yal9j+fWeLcy0OiPevHEC93x2eJFKMnQtZF01heMZBL659XaLGVt3jbf
5Bm/ceJ9SkUg0Yeq+Ws1L1g0husFv5XLlcSjEwgz5SgT2xgycS/r0Xpx6ICtiJBQ
3xiVzQF9IHZbekHBiyThNEE3Vj1o+ke3pPaqe79JoXTIvemtSEsypUABrzQ8N9sk
yYzLuAJD04kah1lxBAkR96/3nf8orkf8XOrkjwFrGbUZv2FtiZYpcIakA9yLQGsm
HfzYgEoCMkBkV4MmFH2OjIyLmwuGBAMnASyEMZ/qrGgxpQkk3R5nZPhixp2hvrhX
pGyM+tEV1B9tl5QmW3Vp7PLpdm0N/k84qZbLNHUQtb6DiDATAH9Byg8nAK5memx9
R0dhE8/6/eqS2V+h0gNlLDXyyCpn33dYRenBArZLKALumKNCXIsTBh+wgNb45D0y
l+gxnDSoR9V3lFm5RbjDP9IgAC5bCBBR60OdZ1yb2o0tCDaEObBmg4UFmFuQXD+X
+j/DH0q7lTGXMjqb+0hIm/jq7wYFcq4n8b1wNjQnfCYuJ188rEu7JT4Q18xFkkwZ
jdCVwTFA0NEqTyemOaadejbH89YiSsrrdAzva+jnm3Raaf9cgvOCBkEr0dmoANN0
c71IaMP+zQFCCYqlnWUfL5zxWwPZPyN8/DQlWuv6dbPuN6/D2LfyfexGEG5hpD+9
wKEdSSLELmGG4W0HcD7n2DTD9Wn7Gd61GnOI2JJP9IJyXhvJThypBDGG0u8hCbbx
tl7Rn66HF62lTfDxe83pqScZIlyB42YUo9PLO1w4yGg8TlRc/DBI5YUyz7U9Ud+3
1h+fQwR+4eACUMRlPEA3YSpcIEWdJxFFsehlej1Ue68qViWIOk6GJbnzX7IT25NS
iok+iG5WPVjFqMNWXEvp5Fb7nbMeU6rO3a9udHT1hlJ228g30nUr8N/xRR1J4gKl
nWN4C2YnQLy7NGrn0L3JoYdjWnvYj7w0dekTietixhAUhj4oc0Hp6N8nDZu4Po3H
m6noNGr/JnuR4Kx+n1y+S8/XO+81YSQ8OCBjw9AwwDkFZcTMCrSuwXBDKfs3uA/z
/c+p/CZJSXz1rUgwu08Uj5q8nLq09WnmkTSg3ATdikcbpmXPo1xtRu0qrMzWOEzW
PMafzDHqX6rw5stSfwf7xCS1cqgQzL1z9VqqV/7ybJxUOzk2iUi7RKvntgU2scOP
z4YZipkGJ7nWttBMYNRXAppdTDLBfomSqWTIia5BKakJNWALw0zwfSjgeorXAwl7
ioP5YQaiXMmUvvGJYYdZ6fpe9+J/+AeUtqK48VdEh32L2Rah3b4wtb5i3PTDkT4U
YYlDpX2w08Nt/LvOxdjIZcdfEvxo9hVYIp0ZUz3ddtcgJl6VGJTDJc6SEvyFOkSQ
hvsG/RNLwOQ7VkrWS9Q2KU90iN8rVuVTWVrrp06eQvTl7q8es/SBoxfaguxmH9+t
WDjhtdylhULQSVC7Nn9pYCSJlhRHyh25TH7vyQK3hgoBFu0eP/1IsflWqdh5k6kV
DxiPsWiFByr9abRl6efhUHY0K5zY/QoRQcSCB1QZfUovRqnvR0Y0HcfhtanpH4dh
WvHmoJBUa1Ea0dEDnJouVsezMjrwZW/mnPVFeErVnqwC97+q88L+PflB+Fog2ha6
HT6PSbPi11DOg8eFkbdotgNaOgUn38IEEz2TjnKoimMh3MPIeJHBYXf8VndGitjv
Rt7GSwf4Uu9WOz9FbvXW3sMkkvOtryYWm9e9dr/siZ3mFJwrVPLRbj5aaafyDj0d
KfEuCnx0YWiYxo7R4lSOVdc3rkmBUJqYHEFBjwqnz/589AgN+IovUt8KV6Em6gXk
Fbdj3HiCxJfeyrsO7YG9CkQ46epM2vykkvPCXt2e2glU6GuD/EQm79v1kCfbE6bd
jZo3dFPbwLe+PF9PkKE+DAuL1WsqA2o5ueNgV673M/PdrplZcA3fY61zxhxOoxei
ounKi/DROposQn9a5CSS1UJ/y0ZDsVxAE/OYCZtQL5tzwPMzDH9aZM7R+d9QBNDm
Tb8BmFp/F7okqyXzXvPLvwi4SE+DX03som+IUH1xkk1zg2Kc7K62AyRdFEaw5ULa
9FYbD7OF34GqW08vdJia6ZMbygWo2GnkB4CMTmUpZxy6GswtVKUFX0zqFX6x/fKF
9fMV4iqib9GMdAfGYDdy3YpcntDmEAH9cUcvbWz+9DrmF8tTCGPQQA8Th2AoFfsc
FSv7Akf3vLpQ3Mx2UiZoDjUO5DHQa34iQ3Yijj64wvjtusx6DQU6gev0FEO3+k2r
McS/rFykymT2yj3h/nmBCHLm2zSh01ZOd4SeA61RbciTvHp0MB8jhpBYFLuH2ltx
LbX3Z22LK19hR0QhiJJFaZhdoSUobSwG/ZDDXEXCB9RHoCS53TajqPquLZHpTmm0
GcRv7YpJtQ1edgpnW0+mNX0DGBYmU2FV6LSxnBwM6OSpz8oshDYUPNmv/ZzMGdfE
mpIOmYavYV90CbGmDjCyUv65iCRA92QPGad6dQgyXM0U/+z3swzDPY3rJDrpeqk2
iZeUuIQcUOSUr+pSeyvGFLYSRMQPDY67yNbnbmVRR4m3UebsEx+ni5L98nHQq+nc
LY4SwedYkRT8nN4cwZv/1fq3PZ+MlooJIqbah/1vN2FWGmSyzEt+Yud763FIxMDX
xlKCrrJHkMYRwgg/npUjCgJ9ZVgw3JOb0Xomm6R189Niv2rJeWWCkzNkBkd9+DrG
PqhdlTzU5sEqEumwvEkPUQziE3m+976btg30pOHSuL9S+uFZY1AEIoPINJLLCZ5O
brqgDc6vzgrsMMBKm8aDYWpfLqb+5KWvAJtwwD+YGwK+4VevTUtLAWA0HjGuGnyn
fC+VQAr85qSMkc2dNMhpPJLivN4eBgnjxvmTA0mKiq7fqScLja6T3jWgT3h28Xa3
HRpONPQYG8qnkMUkemZs3kaGFo1D0TEnN3Lg722+ov1+uePmETtP/hpANqOg4VMF
muGq+d0dv+VpIxb2Rhx/aKtupZUZEX4fJHNi637wxT8ydfBOf+AXw8juUxpjBvnX
Q18xm+kSnj+cBe9OxTA6JjueVS6AFPGadhIgXnjJNvuuj6mVrYtRLqiJ8Plfhb+3
qQO15F4oEUsFbAtq86eJk2/gNqCrk71otwOk97KiUA0NhQ8fobsWnnrtOjHzz/UT
tYmuz9i0icO5ScnuOC6OQlTm3tEPDlbKbQsNjAJpXQEF9XQvb9ilqVeLHhlp5Gk9
3RmXddm1nYy55z/oVO05TNRhuRlZKkn6Nu7zUS3J8rYoYtxU0n+fuPFw/DOn7QHE
ctau1FxqGo7wuzQRcrtbD3iu8yiqbdenriO66uHEkeeGUkthguo8vOM4sbaOkUNG
hvfQGh/xau44NFMWh45B1BVE7X3dS43m+fGzctoUlDPzKsVKN8seQd1qum1aruVt
wXyRFkKBkJ8i0BnTr2lIe02pevn9cw+FXbHg+EIfz++mrM1EhuqanpRpXQxoXaG8
tcGnD9FpCXkXdWaa7L79RPjqeZKTb3VOSVmGnDIQEXws++Fwu8jBR9Kww2sOB2B/
xmVpyxA/+50Jnlr8qmWAPBCcnXkdlGwf6Dv9lKlYc9DDSDcn5AlZ6PJu6J8JUdAO
U0tw3r/gDRCQiQ4eRn9HfFGgn83TwgKMFzCLUd7QDNLGC8p9A6GNbY0KIhn3GNmZ
pu4E9CoSFhzQPOuoACrIJAewIxXIPT5zwjRgsz+j/ppyoI2263daUvvreWTfoVSG
rr08ZoH7zV7EbpH2XOkuAkqqzirqn91aqbs0b+oH6CIADTmLuouUYl+OUrkpkyfV
vuI33a5/sMVdRTj/slAcPN5doJlSvxuqMLQVmQdhArJQffKg80pm+sgwDIMspRxb
lEPda1AuY+e1sih78Qu4KcvnxulKyg+a4XzchIpVFj2bLDtxpKm8oLbv3Wkh5VdX
14Y2i3jJAL+n/iM5t2GYwUuFEuOcoNs8XmTyIhf5KFJpH27A+XI0QgdMC7xsHdse
c888XAPos8S9llaSVWnnMijy8ZDGz3+olX/WieRITkcYWNtBtaRSKvQHH6l9r1Yw
ByperrDNNuGk38KnC8P9dLY3qkaU5wCFwq97g3d/2lHNI+cvSxU/vABrZJwAMCDp
A1W4XMUK+8IJJyN4UajOmdrvw8J97U/OHvOabW5hQHVqSJBqgmRyfTEQNlwOEjmh
Zau3Sm6mHIk+SEoVsjLfirTIgdB3Gc5WtYpMHXN+j+rQwd503qILUtCyC8dZFdRQ
j63wKT1qDBGBcUT183vVfCSsy0vFwPyvikiDj4POHOl72xaSAjHdSwJZSVvpcSYL
t54SI8FTud+Mst03/fO7k/5P8j9CQ2yBwDTHxKPAGwsKacaAefFWILUq0s7NQHdr
vOeJD7EfsOTiEURl2+TvrugqiMln6Yd479SNEt5O32djUXsAnrVLZmxJVljKjVgg
YbiqqsRorpLEcI7JierzUT8qJP2jaZ2Smh/t/XsPIjkP0bPdmHQJ/J0KUeEe99uq
viDqjtL+jn3NerMUuiuxKUkSo0u9BMtQcv/fWCiEt2DegoQ90p96MXIGiSEWnSBr
2qHdOPlCVIVjSe5PbSd++li896Sd3i6LTU5eE5WNK/1cStjVBBhbYAWlNAtZOzVG
SVou54s3mI+V2Ci9XRcFOybpq4EhcEy5uz0k+b9WcMvPoisybIbQczx6/qgn6O4r
YRkzx8oJNKkQinhDrC7zHU0gAk/X/PGAcFB2p38NhpZFAjJkHuxzfrsYpT4apl2L
fGSTjSqJVWBiXNC0GzavhSkFyWgUbJxwC9MpphxzLCMcSCXSSbLYJTgd3FKZrstJ
SQUK+5jVQk9OGt6rwUSJeCuAXupJANWkvA7is9xGqCijB0jZAfittd+q8YoYLYeC
ppUOnai7nb+DjwZMNdduuPhnZQx/WDGVeSAskeVsKrlzitRgmvQL0cRTlCHFiOWe
J5UvsgrnNcIXte5fVhY7beaLHrHuOH41XyGCSEYCoDfZQ2oRLCwl10P2eS5HL3hq
sFcvCSe+tzTdD0W6SDsqZGRrupFo4rM13rOMzuwPAn5EbGGmhB1isjpf7ZdjCqFa
akh6/e3uiI0P1EnMv5cVFp14omWqVTorC3Hru52QTGDG8dl34WPTM4VtZyEb7hDP
+7kN90pck09Ms0Qfcpkyhbzn0jOhickFwNu/QeWBH6KZmbHarGsg9IdOvXErMkpO
nQFIeP3aNVEoeA0q8PvrWR1UIOBMQp+k+ryBLAI9UUX1LgUbXLQ7ssWPMO9Ef/Pt
XtAcLEhnTo8SGMhnhkS/eyfgyLdgzRWc2O1k2GGJRnxiNxVApDytMaefJdgJr52I
oXL2UuHcU1s5IGhwcpgoKf6k0yOOP4jJYW3EZ94KutRMe7KgHW4+SMYwliVT21Lr
GklwNp2Tlj68nDRyJA+XTPqeOZMEf5Pt7YAt6DX690O/T7+yn5cF0hF1Ou2CUUY+
tA1nMJ2GZI8VUOfLZBWWW9lFJnI8qF9K8I5hvhhC2N0Hdyu+ZLY2JNYo2kRCcHcN
rnRbUHmZ8rxmvkkKi+nTfpdeRuQG88hPQ+alpJWPjJlR6EUkog7aFhp4mJ6obIoa
UD9kaf/Dozpca2VH6rLl3FWcO1D6y5pnfd9cWWxthmR/kaxsnBan2LdwX9w72J4k
dLOHO0ESywSDxlEu5l2VNdC1e6tDghjo4Y0lJBipF5mH+CPtocNWM1htCVdkeMlT
fvtLDPyc5OOI5ThTI7iHhAjZq9KG8BbNygJPRJDWUoQkGhIdb/MZ6Zhem2ckgUs0
yUE51zSaLJkqKjNlXuz4Lgs2YApxrMDj0q3kZMV/AEK3nLpDUbI23tlvniTPSrp5
Ct5qNA/W3XSevbkCW7JP0bawMTGBB54W+7FaZTi2e4PisqzGnQ/Kmc4NiBZHSS/e
BjuN92OJwOe+wif3K41IJoaLBsN9X4+SB/mv7iQBOLimtciKdCUVrtbK5wViZqc1
Jh2bcDDxJm/FTYk3mt4ajIgKnrPxuNiIiCh8GxDkMvjKONFxss1wTWgnrlSJ02D4
V+nwHdUN56UvditPw2H75BhVh6U9SOaHTySiOgdEZkFWRJgr8FdsUYuCLLX5ys1X
E7JG0cD+tntcTvXpcRx1B4RIA7GGyg6BJklec6mhlVJ2cvJzrz856m6hh9BPkGL5
lRdCrcSga+G20UxMZ2pEvahMwrGUbd2RhcLSHr46osFDaYO6olpppmkZB+88p3BS
B8286XoLeBRi3wUZw2oyib1/0dLFkc7yIrBiIgKFR7a8qE2KoV9NH8izmNZFZPVo
+mfHGdtwARRQBnG+fQP9nRHRAntjxP8Jif/UYbqMwtSxGRgP4AO2A+cgcFkjyXRO
Xao1UW0y1s1ljR223gqG6xOaUNxpb0upBYE/uv00sSvzq7+aRTDpIEiYwWJf2KlZ
zs+8UXAcgN1jsF06qGw9Y7ZbB92Kd9N2G0vABr1OPkiMAlfR0jFOyVoH854VDX1O
pQ2+wC1MJr3VDsz02cbFMWDuO9pbvwqs4xDC5C3yZxlAmSotZ4gcViNRDRm8fpdA
/TfFRWVnJzHEJQTB755xSPPQ6XLa73gCD2Y+4MKUfcwVb2gpVhThqpBynGF7vD8M
VAiGoIKuD8PnOPsEWwwjqyttfeX8GVIm3Ikm0kxReZQ/TA7LTyxK02+ja4VfYqK6
FqkDYcgkKPHNd8FQzF9SixKpih7NCho7O5LOGKLkxErtUso8uQV737tDC6aIAQ1i
KSxFMUqOTKhwOoAcsfbGLV61yVS/NItnMPhwXYXu9xDt1lnvuGCByDTYWZq6ahpn
ckgkOlxeKa7p6LyO0LuI6d08t35FB+5Tx6VR5ahfvkUTSDqlRoe9ATohhDie0i8f
z9gi1Q6fOIz9HbciKz3foIWhisGf/EPBQWeHa/hQzEdQomGtCFoRtC3awOG/Ebg8
CN42l4txl2FPaGZrhpuvYbPwe/0I57Qru19KT2j/FENFMHHHlalOHkuakmXw+uro
riI7BTwhSv0dc1LSpADsIUieMp7I5DC2qdbcPkGBLMxIj5B+pgks/SFnYVuFvlxL
gGJmyKTcsdpVxwVDBaolacn3GiXxnhLBTgP501U3N91Q9WOBHBkzQrPJj0tDZI+L
jf49eX84ovq0VoJba90Gck8I15Q9eZzxYIUYqdfoGZ7FcfPROLxKsHa4a0ZEuD0Z
/puf6CgwW8bQYzKdQbVMdV5SMItRfeMz/cz9vL69DSDIbBtqg0IovcD4vFuu5aDU
i1yzX13KBSQM26ZecJxp9FxRz0tMQqy/2ryDvuC8VRwg6/graCSUTGOeQ72KjRI1
jeQi+atJxJ8W2HzeM29Bx9x9gX9G69wnxt37w/acCbhbVg7MswdtTvY91SF/5RLR
v9LYy9GOF1YI2Lo+Wc4o+Tzkq3dI3XUmgbh0bEkGD+nnZ1IZygluZwAHPyaSqTAZ
6c89tlUF7adGIBbFlWpNz7jcXozv5bxySq3I+1mkx1ijk6YJdTaE7na78clPKyom
3AR+TZlOYLwXQVKLlWb+lzAPTGlECsnfGruo4t6GoHB6hDCMWVIgbqAjqXUjxNUx
/pfE1o1tC039pGanNvtLLR08+Zv5DySFvjnWOJXj4keVKsSHCmeljwYJlbeqByLi
FrUcuYGnK9unGMMxZSUQUHLv/GlSSGB4ig2pLUeRfhzhMf3dwNIpyC95JijrxlZ4
OKNBQQOsE5Sdo822suNJcq2eI0cJLPJJDeaocVyq8gc61rotPXNwFiLEO+FNgGWK
GPptzuoUhxbos5yzyl1ZsL6rWZP6ZpQI3MG4yW0N1WfTNXgCXUaUW1rimQFoQmXE
3/AAiTd4R8GoYUMK5ZUWDNqa6WZH71pFUleuhhoZMwLyuGNbbrc4kIcM+ooJz9Sb
uwG4u/44JpxGjPpVSYlC3108SIB+Ilex/8JSt1EIEYPf75AQYOGidhz6XnuJloe1
Sxg4R8wR9+8zWp72JvM9IE3rVx7umgfolQ1ljshcFTi0XJ2eJ6YlieoP5/Af7zjc
lslOALkUDLy5JMqdysbpRzmr90SA4jsUg3ZDA0VNX34loW0jF+TtyVQUzg2rT2CK
SObMWutdm09ljqktaiGq/OFMc7U89Mske5soFZen0Vxe7CXAdDXcNeqnR+sCjK9g
r/Hq9tIVUkepCJmE5FCTR5n6z7RYGPw3E/rcS6aHhKa+UKZK1SWluRuTOEKhC5XI
LKZY0HuUt1WS9wzT02aT+DNho9fXBzXFvmp0usS6Gz7GhHeCIMSrdrW6t9t+TbFe
zJKk9IyV6J8TBOXWyWX5O34XUJ4naJ3Y0x+oqi66c3j9PShwAhVn8E6u0Tmhjs2q
WMUXI5RhzkyT1nwsU9JxhZlFLV16dWA1x6ju7jOtYCpa3e/wrF1YQMc8r2ty9om/
h1GEkjc/JXAo1v+TEczU2DCuzeY/iINbuQwWDf1JknpERykH+9qLt6+YL3phAmGX
cb3SsHKB7KHNpULzT5n0PlqsOktEwG/Dg4Tuk2wzUJ4jNfgxYBh0VldATdpd3iq0
aVvS0vaEdUwSK4dEFPduamVYnLqo2TQHYIO6eG4VDzkOlzg7d2Tp/chqgdLyX0Hk
2DidVw4Z84nqkSrCb/Td9LRpqF9Rag/EWcS40iIVNU+zYg3AufjsFE1iPM3L71UP
OtD+khCpwpL/+ld+pjc4m9ouGtq39/3eKX3SaY5iOY4YxaEbFWVQXWV18kR4le4+
h7QbhutgcxvTM68aVbxC4Ldsi24QICpM/jq4kbSM6psd2BPu1BjghI4LSAUeiunX
x8YpWcoB2j8rOFzQA5l242YrBqA9hwp9DIrk/kAGozgiz8tzcFt7OvN1pNBOJ8lT
XRjalwqR0nfHYXRgRqAfUH97m6XbrmcOWKYiUXXuNC4WBNBHC+TXnJygPYcY25RN
D7UH3GPdN6rBQFm4tSVsbuw3KE+HUTBXRAUGshpAK2DQanSOi544mPzgn7u4nT8J
nVjrk6DMgLvP9N45nDfZ7Z6ZlthebyHubB33Hp9hCJWavS6B8keqKmef2Rkpt8pI
BEthO0o7QFGp9va6MZCHRuX3R2t+I9l5yv7PdqWOpjZNKtyPismFqiNF5qenth+2
YtD0c3RhDHz9Sgo9efemzjG4eYuXWBFtLJa8zcDj1sOfQEVpE00bNBjmfew00ylc
iqBiiffOtCE1peHPOw9QlNA8MVL8d5kfozkCmZkfSKqU0FGYnLgXTfazb7DCKFU4
nVzFMrlB7lm1AaDAcWgHYp+lV3rVNvSirH1QvPW+T6XF3OqH0r8DUFSbVXXyWXBf
h8YJ37K70g+bM9O5KEMr5lhCJA6HfPW+V0kdxJllgdaA2HdOy+Njgh53+SYnWteF
FyXDfNJ3fAGgnmKnW9lw3cT5JCtmslkfhOt+AC9d/udQOTwH6NhRyWwYxLorkCe6
91/prRZw22azWnJiMNUXHFpAgs80NutVZF7lw2WyOB/DOef7ReSL2fKcOaDQ3CtJ
SauTpOrZ9T9Bdz4jfHJYJkN/PeAdknYle6JOwqSEmBIAgBMZ1uGPiO5AB2AOx/St
WDwOOWvOgOwOja7vwXmq61j8eO37Z8xueR6jU6f4KKKh9zFQNR1rbXc7U9uGTCWI
yfzPoOkQYvrhynAdaFRaJzm56lL4JNk813MCt8C5KPgYKH7pvgwM+uO1QVxlSbOI
l6jlEs0m4D+uCdUsQ3iBF5bC7YTWMvNovpmYkis+sCacJihyJIXbUjymLtubtcaO
AiSO+vvxOmC3K2US257kmAZsSm9E32xzuhcYEpoD7+DjbX+jR7zy2blf+Z/ZEp31
r64Oq+d4IvMFiCE2NjPUBnc3ruw4wY2OZq1PY/dAlzqcR0oKQvVutE9bw1tjmRdr
vFMO5xRGyHJ/3fbR3eEL7+CdH2vN+eUxdubJ50yNMCDPhhRps4UBR1ugyZSEJEPV
WS0FaWfSVDlabcRhHA8MPy+ir60BDE2oyPekZp+cZG3ypdfb3XuDmHDLgoB6GKLK
jQ7jqOd2yyuF+qF83tfvbC3vmmsz3jbLRGes7PRvj5JREHJLj7HNfVQVrD60Tv73
Jc7MYaEwVEb0zRrra7AasyS0BOqVrgQQWdVtY5P9RoWqJIc4bBLjOeB9HYyDwtEy
zrUdM/0Ycv/rKsOHkzN9mknVSNgKGsaIFmzV0yQnDuWAB/Ak0Q6ayXYF744eJYD4
qiCgCeYWKXPNJrmSoRt+Bqj2rarQr7mT6C8rJQRaUXL/LQkXyPFCBBNgEYlkj3ey
xpuR3KkpDC9n1fBcTwIQc1kSCNwBYvtlPtrOxbmDsTOjTSCsaGzrwJBkQsoGQjqY
RM16hEnKAzJpxjAORIJ27b/jVky4T6Y5ireL3Kggeo6SRERqBmre0sybdIglIJHQ
PvQasYPUGgOL83rpi9TTmAB3FUy1g+5dsT7idUEx9NK2ivEjRnVX4aa3x6dCP03m
eLDMLRsvH6rIlkul7llHNqrtTpu1djMYdldxsxGVFotGH/PKSXgfbwem42wmL8uM
+an2VNK+nxSuh+Iml17yasY+LjBcxsPO1vp5k9fw9Z69TlGGVig7HV0jOcGcHpQy
1H/b+iiTpbQ+CsjABSR7GTxGMTOiU/jalz8FmwMVzTMeDV4htuGAh0PDKWSKwnLV
aZBadyL+LNoEOIziwXWrBxhVPQGjZP3obAwx/lRhD+JxG+G6Y+ihDJ9ytJPbgIty
P6XUxXo3xhp1/+ADvuYSc5W9cp1F6dVPJ6Obuh8Pmxd+v1rzRdrXLAsnHtOq5UAa
hO1NS4oM9NIlNjfegdpvoXbTJeUamF1Oq0YCU1jImoq7qElN68FAy0wACti+Jonx
4AwkhXux2rGAhbf2n7VDLK3jfVhdPST1eGyoZZewVdRcL6m+pTjVhJGjRQPZPMLX
kgfpD+ind9h4GxWE2LuE+wpsfwJcu92QZ8UOZBDFSaGrPQsMbJjxuRNyuTVLugE9
U20wcyEhllIrURK+/ekhT6oTigCE5++air8C4CaVjERJKfIiTX4pG2ZKZKfMgVVv
XcU9YvPNLpclxZwjk9gLMJjbV4zPzZ19LMVWUns1bWR3OGXmvmPn4EYvwWFKgQ9q
YyQD+5nGlpBCTr2RHKgucuHIz72SahBwvjMFjYYDol4NnQ8S0tsqT9Icro8/nVfh
WQUl25tbOcI1FOBnQfqGl8ypHGA9B0ksyjG8yjrZos03+i+NP9LykzvGaW9fVhcS
mGslH56Yux6WAuw9fhpqfg6lTS+AVW7sMof1SMki9T85IoQjlz5NjikIwwYaYcRW
eHlkDBF/8wFlnHDPnmd9FhqdlnIttLEvSQASqVAca5cTl5nvDZ1HjuKhhNrjmuVA
bz9xA/KxNTkwM0cCdqlWlC3d5OK7vKAjK6J3cYtAUUp9OE5pEwK1CQiFoc/FKb0D
LyOyB2KeqPdLb+DhNSggxNsUNXNTavfsurxjCTNYJs5JeIN+xUi9RYQCEJNW9ugs
pP2RrF8GH/PFJAAtgnlIZasj4FY7KWT2y6WpkpD5QD1JBgD66bbaFnyjZGqm8Q26
n6KHRENprrFD7tGOp/RLj1r0xUO8uBzZTd+jUBzruQ/4HQq78UF0DztEB/WxgnGo
GBjZuHdXyuk1QNbyZVpoMHD0l0iaR7cJclAOz9RleMlBRQc4LizyQANweRXANtG4
UjPXEIsN381q0jylksFvmB6M+wfggXPtTY07VSy5cgiM50fag1XqkrY2HTFpTFJd
RhJaVF+9e0772LbYW45DGIonqUdZa2vDnqUSaXbgFpc4xbpfAPmUNX4oOt/wjoBe
CQ7xGymIVzsc+JZ/y1FJQDaPwf1GvDwTt0HYW0oq/n9DnRu4HM1/bMvTDKWQCfS2
BdpStBGsXrtHThGywvrW/2St6XktYjdm15ajaCEiWFT6YH5hv5aBy3fFE46RpW+9
BPIXyt7Lr8k/Z5hV2ou1CuhuoLIyj+Ec+FHH8Y9KXuPo4f+26wbfHvAVIA4Uxd/W
REresBaDmk97Z6xNlxez1rOPhTtLRVUlgezScRuXsm5C8uTMpmF89pWT1tlaps2N
+W27tIPg2jYsQkYLjuuXaJ7oNX3Z/R11exytmm1KGUn+eKIXVugq6GGVE/fQYcez
Ihi5SCwfV3JE/AnR2KeBxWdq3rdwmDbyxvVIc1JGpxaM+pnuOXLrPfmsb4AIy/w8
35zzfOMFJTS6XD/QWvVcU25OUau/d9iepLOtA13GaM/wjGgnw/KTUNCuNKAkgvlb
vpNXMln5N5AjC9VkFhuO8YGPoS6KZSg685PImjF/SDDo1nEUasRGwoWWfKGKn52Z
aQoSyoS8ApSm2l86soLHVzP+nLzfU0aj52yzeVVKnAstN3pZ4WcfrLRQL9fJlsxY
/KiRwx9T0ck/44FOlswrijAgiatTDdY/26wny/aseHHWgGXsQ+gfAY4VkNYfwHST
HF8CeILqWrVarlDKUR3SZBVuGn23bky4bEUAPiYFkyleh0+IUka4syvXTre0WUwR
DsCvsogjoz6ybtHSSZO+pm0BUC1GS1GTlbToafNXcil/LgVwRxc3E2ZaQmbXIOQN
UmdSqGYw5R+wrOaEusMCIMjyHI+QPqzdG0B6LrGcM9l63ouNW1/5uk5voTfV7/C2
czpzmAAWJAuyJhqqxxOmPw3Z9jO8RT0IEXpBVF/dpIZUYrgX4kuDS9GjQrWOjsUu
NEw8N5OdBTJOzCns2Iyk86t0q1D5102TZYwCL/XP88xSXi+kAtUjbg9TzDcY5ECg
I2qo/IeMN4uz3U2CCRhQ9fumAm5VKbRBBG0F0XXRN6j1Y4iXLOZmL/8pgr/Ql/f8
IUC/A5ZD+ZFQTp49Pbpg98JB1xX3SHD4G6Ri69Ex11Jo7ncfC5CT45nxWXWVvUPu
9oU8UE8InpyRfUgBemSzRHuWm+hcglJNTslRrZLftmR8O/G8AinrTe2+ER3mbmz1
GVjKJawKutcLfnvRC7bGoOtKxI8MIlHDVi385qeD1OV1kStUGnek5D5d0uxB0RYC
WrAjYR+dKB2QpnJ9FrezwajcPDbIqVC2PS0F4GyuIlS0xctixafiXQEfZUoowBjZ
Kd0jFGw6cjl0XLrbK9fm3dzGuk01ZDYrB7IokUVZITykMQT9NwcZxa0Do//tHeao
VlMc3P2CJeUZZe+WjJx2hHC7v4zxcRNpCso2hF9XksIDnDtLlqgVxsGBPolsjD8Q
DCpSM1faj/y6cjKLCUIHNPr9mldTQfy/OhPCSkZ1kV1Nza1g3WQJFUvXO+yqigZy
THI/I/RRWwKsyZbli/N0Se4AR3AFewsCge84Tgb8cyjHUJ/NZqWAHlhNFHkMoOF3
23MuWGMRKm1wAueDeDC9pbj9d5PNaJ3KEYss9CIacpndP+YA6JbmdxF+PZDvHtNL
M55Pj/MNl6sg7RfHBl7nYVsIV/TdfFYEZeR27W88pvKNhM5quFkJPXKh1jhtUjq9
hD/VUBgePfOotWvtkovRyTwpRXtIgBmQGlnfmUd5mY+xBkdUBqa9PF4qDI7++URk
l1+dHA+ipbETXW/NBAHcxDO7TKaaXoRQy4FkkYmyJxdolQFD1Cc+/8/5o2kODvTE
QPsAFtQpMy9XLKgdNzWFQqfnwIlbcVRAshCFL34IhSGU8JuyYn7cESvdSo9KayNs
wm88fsdOPJP/LrvWi+OfOUG/zjlSEvulcnMmPzpU3tIFz1W19dOKHGoYf2rQ92AB
wjaTaX0Ipmbr4lyrLCnOvYaNhM0h2dqtUX4BrLWVwwFlRDYumqJ/EBk3tathqjo8
uns0Woiyu4h0fjjadwX4BLmzWauzEY3cM6iZ4ksSqbSgXFnx7sRoGf80OTJiGrjI
AW0sriSAhe74B6Rnhi9T434YOJtki31rjn8A1yvAYW6HQwZEU3IX2+1QnjpF6SUC
wIPgVAjs6+DA6YLLpL5IxllI6kYG90M2J/tGwFSBBYAhgYlyRbREBdw7myNVBBRa
4kBxkJvBz1V5xtbAl0OAx3YP3aKhBXEj4UNUX+5mdCbOZf9i1OYlqlXpF1pRRbZN
GY6sY+DvGV9+TuyI+I6Dyj6/EuHiwM2VIKeB0osKUuvAS3EW5Fi3dNnPRVxOXhDQ
WLn5z+wIdGBzEhmVilFC5hiMiAKH4zrd1JCnH/4ErB0E9GOl2lxtiv4n82gpy1g2
dEcDrG/OyPhmzH+9En9VseWi627t0rok/4YFI4Kb+cBm8fTkdUQ0iV213SxBxVqi
XNm2HrdrkWWQ8erpZLgDHJGuMR9MohUxT0iH6cFiRWiG6pKIcVOB++GIQK+8Rrnu
49sV0Io5rfjH1Z1nCt4nN5fougwrl2VndCMqIrKaO/mWyM3TslKo6RtIn2OziGvG
/ed8dnaH/R+hABDuGK9U2Tg+THFXpXp4KhMUe3QI7hmGbGjsKybDgHLyM3P2UrMw
rqWqF2GGHv5QmTI7EL5aS3vs+crjJ588OM4I4vDmUiELvvUrDB1sF/Hza+wFj1Wn
DK4eE6rn5KAjEbwztzvpLb6pIHz6Mcds/K/tzE2ylY/wtSpE/1uNX/CYROOP8C1e
+siVQD9cPTiDCJHvqvUFc5e4ObExyO2DI02AiBiOmXiC8lrsKaok1WYEkrwmtHlE
cB2FWO/jSmFdPxnB5/O7nAIFuNmSvSmaQ/8DRblf34JuQBuic9o/HWNrGL94bFeN
BL/APJXpBlvRLrqom8QwbzeqybOv1kgkMozJEtSh7PBDugNr0LCgFblgFTgjGRrI
EbNhkNxypldQYX4tHP21lNJwJJLGkqChmgVcgFmIkUHjSWaYCVkXToIIAEPgQTyM
VTm3AmoVlA2mTeAyxjAQaslINwaqaA6BU4LnH+fc7R8HYygvHaw1wJ64JzFhw/3D
5Z8UZTCEHRomqJ5JMcbPFlAKttUQ4M2KCmLivBYKmKqLfWMQ62E9H4XX1sceeoRb
lQrs6cV3ERDhOHkMqbGin0fxKobrCIATSneJQWRWNaRLFutjQdTKWrx8fQgJwx8h
lHnSQuJWw0JnRjrjMi5xG4a71Q5TBEfd8StxZDUGAurYOlfmmI7fQ1g0e8p63A/b
u8no+jqCNkqzI52vNLw6I4rhTDQ55SArQhnkb3GDtXUK44rvLGDF6DQroLZ0Bbxg
RmZOcjYJQ1f3KZuTUZzl09VeQ0Ot2Fq3xkfchGO6EvQqVimZJKI5IFajZeJf+18f
cQA97wdqNeLLG6QY95bOPuikKzMjaQ4+J4vz3/CQrXRbK/1z4KGpuEt2eYlTmOiM
u1VFttvfa0MvOIISaJ6aNqVsd65gq9OZQE02dQFAhP80ZvStwdif9Vb/+1ncImB9
kzt+uzEBvDccuil6FUBj5g8moFa1L+cFe2ixzFKa+ysD5R6W+fzR+n5vLCQ76viN
trSFbYV8mC+6IZGvj2GcRx3SZTsuT3JouxfvB8pJvEWqcAn5mrgOa64ZgTVsbUEk
HEymxMMdutZ6lKoKAoViG6IuFmMLpYgehh5QqjfYj3jwhmwaDR9lQUhRERIVmnXI
boTZS7i7zt62p4vJ35ro0ho9zrTUO3oXRCDJRGHZRHpP9emq7iCJdIo4YDnmJCGY
TXMIhrrDq0Q1eDHI1yAoZTgP6cI5pJgPTtZHgstEJmHTWBTlUu+8xUF7Wb+n5+5H
uxS3cWLzAgrshrDs0WeqDHFFyJseIW2UDqT1ZHDwdnBaCed8uLAufKGhBhLJdEXh
8yTJqZtjNPEDNwmAFnWs2Lff8t40wsvTobBr5ge0mt5YkAnpNer0S6KTsM/HnMYC
jgBvoxmZ+/C66HwLkz8HUZiWVVfaft2YbyuLvtfmoneregXF4ZZDNdgkeLmA9Wrn
ogAGh1ELPYtsk5w24OUjcBH7tU6WPw/fi+w0vwAfy9fzFfBd6F6YYOEphsmd6TaO
yyTY6fjwXpgJDKzvT6cygQ+QWA06Q3ig9xnP/a8XgDIoyC0/x0knm5yuDUd7JJFE
BSxATI5Ki28bZdMKPUBIrlDZ5ZvjCQ2AgfwZrToPADEFVaKpDE0dGIbUCJKEtPdD
h4YB50Bdv7Qu8IhuRvChB/aHF1IpOocxWwm3ZjO/b4QIRsXT8VH60Q2qtZT4g3g2
09ld5ggIvPuXYWeOqxGGdFobtZwgsiZ420kQfyAS1gIwFSe8hlZSDwKPz8K0fF+m
FY54xjaXLwqTcaq1CoEF5R64QQlrOz4VJxJwa1n0EYNYKzKe2Vgk0WPZrUThtbaO
tpezLXqmOZfgX0/dnAZ0JL+1HUuJKvXB1BzEjk5pSz4ucTlDxwElmGZCGRYNPQKp
M2HUsWPScaNTP+vCDBJnuUr8+Z0PYqLJAJkPvDr+KPwkx/OpHrkPpXOS65hlpu/u
CeUeJpWw8Cf/FdptQKl36lcbrizgQnHe138SQbpVx1a77ONTpFUARim9XDAMwePL
5hQrSm3vhIjSwe18q81DpSRN7+H8yU3Hmf7l2TDueJVuPmhgVkrV7DCWD/UvrMZG
xQn3HjzfCbUl3foJSXyNdZasB2lE1gD20qCC+5ZZqqB1eokZKfWdwmhC8iKzWGEv
EVplsAMLfKk4YrSNyFPhyhYGuk63awCNfOD09QwoudOoOJQgFEQsDoGyDxsw099a
Fwjn50XtaUaMu7+t/+A+9qeanBnGBTzl/xKJxmWL92A4keoWtGPwu2TvG+s0Tlf0
f6eSmxJeUqbXgKyDABgWD0N+Q5s3McGl3QaOdLikOeu3R/CkaIMlZMslZQ3lFeL9
Zr2qf3BNqAlsxCYJU9ytrPXkNMGGaT43Gw1CU9OWiwhAPelQruTv4SbKyI2DEluI
H6/pH6rN4Bv6jmMvuuABqwkMPhKgwz3dqgeQZR6ZcUOgaWzJbkEeX3xkuJH5YHy6
O/k+zB3WZ0uPCoXEjLEbkWjCWi2WcZS1gPGj+V54Bq/XQ3g+1ZT9fTF8SL9HpK3v
oCN1kZZc0JjYq/MurcGsmckOosSwYBHoO9Dprx+zWKZIdFsw7pjzP/JdEgm34Ajl
5PjdqJv3oBOQxPmkzdi6xROPs4NZhvdZDKJtjX6JC2c1SCiwkDTCiJYKVT9O9oir
nQfUOEmzGDiLuPYHNM1QT8iEZEtUkGxsP5lcQ/htdYuKqC9huONUtflvi1Tb8vG1
6rubkA0ybrgu2c8T8FtM9PFZamGOE+9l22sC5PWhsj2SSp/gVgqRCdXGA7QovyL8
yZ4WmxmjqBAHWAldFiqiUodTt6CWpoKNzgtzVlxwLap04cKP4GUDEgbIiBxoOGlo
p97s6JyphgClJjsgbHhU5XiAPyyAM44coMe6WwqfKO1jD3IuAS4MKEBdgD2saiLi
Wt9hyCBh6+mJuDwxQQ9mCyt4fQw4YcPbW7kV6PVYIEJA3K/K9BgpNRFdytbEwyWx
0PWcdIUz37k02T8Na0oESxiGKpeSZXUQdPbOiPR+RXrgJaEa8PctOWF8RPCBWAf4
mX6TMVYYp0sDokRTYGLq/zvYNzbxBIeMjcoFFS01d9lSqeCalkt3Yud8G19sX5OY
NXLLyETpeGDZgFABg32/JNKTTAIsKXW/SOIx6cTnzsc4tySOppXHRRsa11J5gZND
Aa1/UQtP/AGVUV7XGkeV57ME0nsCfMhsk6dHlINokwvZQdDrOXEzx2R+eKj0SSuL
56hw6+uuRVN9uvCPY+51/9Bx8ImABVGv4VQLu9nSWADSbK+WS10oXVJio/DdEdy6
baic8olQxDIlVcTMSvdDi0cPv7WdmlTnku6sha2S68I6QzuVB9DBX2MVB0pXqOAv
c51KxxNIynLPnuL+iSXQ78+sxMq6c7eMsPnMaIyN8bnsmEZuzutuoRhNmkBoMow7
yqpJS5CbYMtBIoFtH32E5du0/6yGJ3r7MK6fkPA7OHOltzq0/BCWhIUbZizCsQfn
PsnoN+AHko2WYrlFRPwnZt5EuHrJE1IX1VbKGigC2YbMCs9wSwVyUexHakrE64ki
KWFZbXHKgQJUo2Nwe0THShqo/f5EJpp86jDwacoaFpOa4J9WwsE2d6mnpdBjh0te
C7J386UEY69+kHj4ZJ284jxLuYjxdnXMKjB6N/M2xzif1AjntwxMtgjxx4jayt+o
bycFch7GCAVyGwa0eH1IWmGHNE6/2T7lzfhdCEgK48ufdQnp+b870LctNW2CXhGs
0Q6fgYR29lHgcOEIJGCvwYsQ/QSjrE37yNG4VXDCQO0rJH9t4WMTLrjYg1ZsWaAx
7QnSIGiDvD/ffVeMnK8ZeB+1oHiMo0GemvHxC5LEoPRBj5LTDHPbSjLOJO1x+dWi
nJ5jtLt1soTz1Y1sC1x8Qi15DAosvhfoys4XBY32boHfZ2FbJ5QGGwFtycxPSDGe
0Q4lvFG0WIUkVu9hIW5bN7fTO11rjwjOZGTyHTm+dmHwwo/lggu3RcN9XXrCL0bv
8ONqDfImkwtNLHsDOgYWXAlxU7cxwuKEnT/tJBp5U9g0v8dRHYdl7qhvT9BesZ5y
2kraZgYZyr+b6LCLOEtvbGYGXl4isvCsiTLGZhePBojL7jADjSlnPa/QnJdX3p3C
egs6L+ygSzgp1yg/gxi6cOwRrU+rzeINL6DmHc7bPoiJ1TWqZUrpqnpgnGVK+K2Q
BR5id9uKLxm7ZJSiErz9DMndyCObXAfMrXceTEs8ssHKyKlVGkFAoiHQ5e+SJV+I
LDAqVgPUs2/EplBYvHogDmPNS9Hi2EQEpCQAR4lsjKBIPDCuNW5PNkG4/NIo8hVv
g6CiDUb59moo1/kugRGTXrUH7fOUrIO2UmOvFF7DL2ImC29Wh2lurKj2ulawT5jh
mDN1Esru2tnV9uBVSoB7RozGJGwyy8L2ElEcTrZYc2Yl1eqxVSkJwwaWpqVbEmEm
jfWnqdyQc3a3SsH1AliZz4STZBdbTR1ho59rvL67jzqPXvpLjec00kEZdQgdcatq
ER0uq1fWhLJInE6QmRXfhH5Pd09sPYtJLaOx7bIJQiePUia6+6YkuJBk7b90QkW7
FqyZKkTrXNlDhfPc84YHlixVL6mRC869Y3wCIQTP/KHR4sTE0zTo06HhQ1mNHCom
nFuTlHNPTaEpSFU4LJBgmIhDx5lCNiKdQK9UZIB+h9YdtBEp7UngoPKGaqCCfBGb
ohcG5R4dBIKhsk6ugEvdEpFDD3o5VRLC64SFW4PtINpg+pEKpZCVC1NzIvhQsEyt
EMczHYyIXKryUAXQVq8DoZQCD4bOncre9Q4dNrwhVeDIwDhUNGVp4PEpyWAC5H7X
rG6mXNF1CpP+09zHBqB5fFefJuAO87G7hbt6jCQYhCMbhedj1cKlOBTc0p4kBOho
NT5Cp5fTM1IG0R8TdR82RxFcVVBUQ2nOCDeCIt0w1qA3qWPzHdzk6eIc3V/28yRc
Gi5pkb1MrLfQD5Zgrg91qQUUYHTwclgByMEzHdTlILTNNzmBw9q7IA4fXP/wsHcI
I1jZ5+Citv1Ih6KYB4hn3HV8ZSuIA+FdIoM7VAYdmhe4FjD/I2eDmP7PW+F1Ey9A
WNAbB5mSfZZbaSxvH42i1t84wZZSFs/2JNBWhKK6eZCj8obeOS9TmZQCLKArdyDK
YXsu20GEAN6gDSTpCibp73noJQpZ8SdE+hMHi+ai9qzm0dvCaC4DrNEbQwdc1sZO
vpGBSMbLGx3gBAXohDRNp9k/qETR5m5b5GDzRwRu2Npi4SNfL9g4F2hONf2aRt/5
l5SRSeMbF1lEKkePIbnI9g5dRtR+u4GXATKa6tF/I5uHJGiF1iOrdq9+A58hxUYr
ioVm10yokbeYJTl0Bo3wB1rSweZl0RmDl3jSHA2+KnD74EIpbKtv6ONtpdtUbz6F
dcTr6dq/upAnKcevk559OnHYPsjP34qpBvHga1ZDJF8gm7qOdyqILMnrWH0aBD5f
sSWFkoQWStH1nrcnlKrMhnJl/DH5X5l/tI2vKbSUsut0Dzl81yRUHwe+jq6Qt3HX
FMODZRqocBsQJqEyrX/D1oIz1Sx/ThMw0ZyhOskXdyb6qUXc8+Yo1Jajt6exm7y0
ZDP+NUkI5FzRzdnr3JjNvwAzWsTWrCz5wQIPZ7+7Wilw2stf8tqnKZ/iCZl1056/
Pb7TnHVHyelYnvhYRzxnJUa+2ksA0qxFD8Y95YG4dv0kxc8Arlhipy5K0/U5bb+Y
e1dpY2PX36uagB6/OhSfAb3enNqLVh/1mnYqJvQ9UCAPQ8Ix4sd8K9yIC1I8CDNS
1dmTX3jTYA6IyXp+UJJdkxLla95OgTftu31e5TgpRPE3E0zz0ZtFzNVRWLnlZkyk
0r/84JWpDx59d+t/hg0F1yDOS8Tjrz8srE/GMvFQtohRp1JNAJQVRDiVwCEBqp0s
jfYpR9Rp2CIb09VlBbxP/OJGsQkdj5yEDuZ2FXB+dMQ7TAfPyCvqOKFmav4Lgiat
Y92IX2z1ECKVnQXwQNuHEHAAfHFYfhE9ShYCXMYGmL0f8A+7NEO0jMTgZiDYcwby
YuDcf92UaV36iIMyN8YnAg9YtWCoYc43e1x8MSp4+bM/uEVwNn8MlTdekSM8tT/d
dSmQKjg7ADSKY5+xMqQD5yJ66x4qvIlkRzDmPTJ1Rwqq2M0RD3MpuQVAb8DejVjU
+G1Q4wuynr3jRFU2KSdfFFXL26p0jbp4+sU6IyWr5VGLI3kPVYgXOscym1ddiStB
AWNn4pxcb2/Z6lUZK4OBRCNUKla6xpIQ5LiWgajUinrPvlIBLz4gHAOjreF3+QFh
wbT2721j02jEEnNgkmZU0XmNNJWUaq56WBsRRPgeBzKvzRsyUtOnR+UaKCe8baGF
AFwz2I4EPdB/5fuOZt5Fr9shBSFm66Cy82nwtmLx3H3pRQoXlG96GbMwn8xelkSb
tAFbmyR75HC1NYNsqZFI6Noy9lkZM4UwPgY/DtZOwr/DxRxmi05boQHIWgPLjUZz
B/RAuRGcmO5cha4PuAsG5+pWxlo9CDo8xWtbcgVVG7oasG4HsvmSuW94greieEWe
mP+Pm0NS1VxMPWn4YXGGrHIULop/CkUPCu9geQF3qWsbHlrPVu6ZcRUubUEhqTFy
rwMJ6Fpi+eKyRh1W5A0+MpVk8EFs0fFYxqLKI62IuUkQmuTCSCF/mqPFzF8FDcwc
FCtiT0YP81xMaW67EbAJ/OeIcvuGRugMBNoa4iWd3bJZTT8XvRLfecvvl5NKZ1ML
Rt2L92+uL+bvTsZ0Tq2ejmZ+23+a96HomVDTWqDZ/7+QE2IoDPaS9tB28fr6yuT5
97Jg2583vtzY+xRH8qtZ9+XSZBW/bd1syEw5GYfbOsiOil8rTvLPRoHitoLwMEsx
5e4Gy55VEYU67Io0ubKy9fvhd/kY62fCDeugUQuoVsQ52ZSn6NCi+9i/B7f915iC
4boh7pgIPPT2JqmMknMlvf5OoWuTHuNPc9DKMUVlMdGdduu3hxvotPzfOFird4qh
OPd87wgSp9Nw3XwVLk0LvePAsgjTlxQpYgpLv9Z3QQow1JExSAs3cFLQI0V4h2yY
AL79uCOpQl3cb+WB2hxdvz40pZ6WThQjBODH/zA058WOrCmKDYyvW9sMJTWwukX6
8/vKZRWgA16jEDZntc4cLBNPvKSTLS7NCaGydvPIZmHjLDx/ufwyz4H0kULyhGeo
aQVnKIgkaNleIQArGz/cY9WX+W0yrRGXnQVCOuwOllc9BPTCHfTcICiPYoAtDdAb
GMzWxrWtxXVoz9HULZhtEPk9atDgslGFg7EvaNYLwKKrat1SxxsMJPp8LrZdvZoR
Jih2+0Qd5I05XuyO2PNpEnMT3kfKT4iUGma0FIVi/ptnhlCkfonY8/oxo3QzFtbx
m6/TIEd0EXix7D3OCKnI4+lPDn/qL5YvC7wPXGc0D53jnP9WmZkntroqdPOfm7xX
FcI7PQfht+UItThkKDp6ENWb3wL9QlDuMRslGt4n0nNFRVQ8oa0L1ejYIxN62G22
hWcUVfDK+PsSvkHWJycTqi2s3/eHw0KWTAaocpLEIz4yrmJbBjBJB71HsMaLBo79
mZZwV2XawIijHIIIrYsMGbFaPmDTp3h/yTFiGp2Y4Xg+W1dOGkDFD8h0YdiReteZ
M4zonYmtt9jwkQTume6HzRTOrUj52YSfjUb6I5tJlQ5Y0J0YyGyQYPcrYdSx1MYJ
hIaxbCwwMbzKwFNIvTRnHlbkSFmocyjUOyLgbT9KJJuTEh6TShtnd7Qj8WLYQJ6N
/uZOsAt9oF64TD4qeHmKWIjCaSMXC1WEZ5lsBfiiPgkVZGYn7wWOjX0pSnTR0EaJ
dAO9t5ez1PapGLipoZTFrcdULzwCY/9FQpbwEYZakkHO6SylQPnXD84y4ew9vfeQ
Fc5ygUBiyW7zSwCk7U2E+zC8GW4hMusM4XqfSwvi1ZzbppIsC5mY3tNgfsOeVyq5
SLG+ZDf3ceEyQ8rmLrN1wXgt8FQZAaTrZnApWGK/N8tA4aFvZ9jgMaYLIN0OF0rH
Rkb1U5qE2+oawn5zFJDN+FLPd03f5XiWB+PgEs+mbBQqfbz8PPbTXcU+SJ7gYd6w
/4atNcGcJpO8U5cBSUXv0BIjBeIIgdvXJNj3Rop3Ic5Tsf2Z9EoXm5CaRp4SNgfB
eLOCFoMk4Az7i+ORBEzL2nfHzSGAlir1Z+MITAdrH4oMk93vfeqLCG02VFwbfLEs
DmtD3dRtqURMoyO4bzGFJC5RKuEEgejVVfIulvzY/3D++E5rKJ0QjVywrMkjqNk9
9YhgiZxVFYYAA+162hwZex6QUZnvEEN6AwwpsInCTXA5Rn8s8DHXv5wypvIVwugf
Nb9ZJK9lT1GNJ0fxrRXCNE2z4FPZ7CczkwkCXGcrAGtsqni+uF/CooqYq5XsSl/h
Bbb4OiihJQ4fjIM0M/7CVlj3kYTYLWIHLMELbuvukdQgslER3HCTim4SdE+4kMFx
tfUQMF2izs2b1rkHmmWBDFsK1f7PeW2LGA/rwcZtQyHo471kzJmimeEE/sgR6G1y
w5QRsl3csqpoFbGhJOE4+HN1LRLcIPiLJgmOFWbUNOvf7bYraeAkEZTpr85tdD0L
iaKxQYnqiU3Hp0YH0ZfE+poAopXkO7NosUko5L87WJSnFrtInXmJr07B4FDZ9lxZ
mcDz4WhW5hfS6ZNK3GXR8/6OX4Fft5RVhiUXemIJwYi57jL+edUa1+XllYwL0AiR
zLxWZ+0ntCOrdefRuFzPlxS8ZC2OcCA9Vc/2Cj+bo+3ZPZamcL4nAZ3ZZxcXORv6
4kXvPQt9Ol1e2w7kTwFLg8FQjzQZ5sQxjk0dtNbrfXKlYHGjQlcdasFECTUFqqGp
bM+53qd5Oo0DfNhYZMac5cIbSQBnpn9c+a/U3m2B6v3TH6Dc5AV0rx0ywfSRAFdK
b88W/btBj4VBXKHdpZyj6Qk43hVY/T4junlAj8YXpsBeZEXc8VwZso1XVU7bdBrt
Q4gz2yAs/HrBrY32QspFE1y6wLOuYfBqjpLNIYIQ2/c8nilBFxMqqdZGGz9muoiZ
IIL8mrwufiy0WO5Adhvy9AFHQnw5DVwRzzWSR3/q9yH+73eQgEu/w6Y+SBOsVHiF
P/id7brMV3KNFqswYifECR5Rr7+NEO2sT4jfWDL1fUpZtHPF9DhSyw/HL2CM5Kta
CFrtbe2aJ8k70XYm/3tH0+viJQEmMHcL4CtkGUGCpRsDwqTyEinpKGubgXIeA6kI
yHvWltuVQzCa6RZMHIDIkWRPffDkuZH3ERgGgCR89ttNsnW74HLxpKWnmk5lq+4k
0PtXs6TKqOmYuwk6+QDsBO7xndIVF4zGkWL1MoJB4/b9ZGQC3esj1OIxtGb6a/M+
U0IKHw+hJz3WNLyrMVcFDaWhdpn2+V9hfWKmZJ1RKl0N1Ohn4QV2KluXMI1dqcQq
shDp9Gkn6UMQXNZhT6rfuXj7j8QqdKzzFGdrcTad2+mod2FtVRwdB513WVxz7TZ6
Ac+tqa8NNS2JZrTHK0rHoU6Z6g6nCRW7gtV4Bdwpsl6jb4ogXj1cG/zatoo0j4xN
RSkj0aZWqMqCNdw9phGBwfWbDCX5iRyWqBDmdELS4WULw6b84VXOVWi3sAK6vwlO
hD5CHgGGrrAaJX/Ewl2qxhFT5xNFVghkwRqcfjHEMoFVcrnnjyS+KjrQ+iD1SUZ9
N/x9GgQIneXX78XEJctZiNJXcCeCOJ0aHOLMAFm95hiCDsUUjy1ZE9mMb6skdr+q
wx0uH3pV3IXOkfTlUDtqhPqjtGZnmS3rgPyblpqBF6cc6VWuVTt+QuH0UzoSUvfH
2vL5BlRoeUgWj7QIlptZ3WDMuRcLYGl675FBk7eTiJFf4f9lZnwQmc67UfB83txz
TsN2qVGzdtu4oxVYKqh+IL4Fa3kICaY4w2fEOeQJleEb9RR8USit92FZjEGFih6c
q73Nl4I8yPJCoPsk/eqwQ8l6RSso4Q/sz5yuFQhn4D3ZEXloy+I9Fmm6xi77xHw/
UCwFpgWchAtCiNgDv6xxgfao4t3vfVRH97ytkL/Es4eq8909s94GAgRRE0jBTFMB
e94GLjkjcqjEjX3rR7JPgzBYF9lS//85zv3KrH9U+Xe9weFcljXNZvfVH+iyuXYy
iLIUtqgFSGJTU9WadFnxzRxayCqewci2ITwxUDtXJFGHgIlKRSkMAv+Q0Qq+mBwv
AoPM59/oUrNMLxDlphN9rEDW2+aiF/soUg289J7fHDxaPU6PclqyM6yBhhMtXWyr
2zcgjlXoj7gqeItxa5TxAH2IgbL3rRE+/RVfNeUBTs+evhVn4T8zshRAC70JpIz+
1Vi0KVe2fvc6OZ1WxLsX04sKf3h5MQK3dxANSxrMdQiA+egIEMdzeAwffckZVBJW
lfBjJQRjzoFqB/T4TvrKiaPGBWaj/9vPeOv0aLMpPooAyjIrbRAS8qbLUKmMpMlW
VpzoIooIC1K1wtvEKEwn6pKajJSBXnDUkoRLfTQjzFK5RwICHipUxKGyPjjINeRB
CEPCLyGiwW6WbWxtlqBQhvb9B0LmsrJn0Lovo1WpOBdf+i+TrbJe73tev72Z0ytn
biFc4t2oaIH1W+Td8nElGLSKT80+FybGJu2u/9vfqoHiafTeUUQ07/EYpSMiKW5G
tUuqOppVtn6YOsJc0JP119fJAIdflgbTDKhdR1MN1jR/eTvrQxm5SeisluiYIKLW
gpPY6Fz5NHk+pf3Xrop+PQSf6xiP3tcwl0vq2x/uD/4mh4wKyl84ICyQHn4u7fsH
tbMuTLPAIPw83W2SMOT7VbL0evWTFqmMvhrMPHhxA1rbZJudpZNhESx/naMvl3L5
I1hHKwiBYRZda1QDjbx4mpGrHCDVIRUXSx3LQPsRS0HD6OjRvzUBpmuvIqwbcdLL
bKpIfRWQt7znHvDCbtHWEQOiI7fpNvqn8GnqTvhsaom5vp+SMRzjDOnzlSU9RVAY
unaVO5Hbzu8bzzn97iKWYmyfbn3/QybfLVnSYbWGMMduS4sh2URzmEpm84lyhAxT
ywh4l0Q//K9SJOtJb91wKp3pCAOTugpLuLK+kXN8BxMh1RXkVLQM0EhoviDza7Mo
FejLNhAWYwT9cft2NjWPrRjf0mCBf19mNRkYRzvl9K1l7t70VwvoOdyZMYM4rBZF
OlBGlnRTV5L4lVNXfH4Q7r42UGWPshTREgmrOnHQksgGsX1fBM7dmw4cE/OOMZ2p
WNT2uMbylWp3lx5v1kgSsrAiLsSXIvM0p/Vt9kKnMpYbRdnXxuVMagshAoXqf/Bv
Xrjx5dWd1HS5iA9Ly8hH/5RS1Bunf41BKWwnkucSBSnQ+ROCBn+6hQePXKU0hbI2
fvsVUly0R/YpXUGN07NMCK2z0IHDTMBh/UtrsygbD9AiPMdC9va4vIMAD/zoBaGV
8zn23yvBqS3LLCzOgTtsS5CTpdxe9xrLaoSj5ZWekZvs8T9tB7xEHme/AujSdfJk
9scdULPP9rZwTfoS0Eb+x5WXIohcmVtIDGb7hOqJTXknvHFCBpxpflQ+DU1kSQx6
7ruq1ACbrb6XprfSlgtiFIrBpkX5UjnOb09ZufUAPKyKz+3hTRPy5sPHrgw0o4sE
JmdslEtka0BX6Eis4rLEZItmIjO/lODfg+wPYNhV+wVIqXgYUOfB0pvvxTL3vNbU
vT8UFZxoAD0UqHPTTvVXcQtR038jATJfHk8UCFaE3UzxLORAWI/o8z+oyOON+O1A
BOGUgZY4WqAEo1PID4ojPv0C3wNHAefUuijU8ahw8FFQv1borrkbNVU/7bn3Y/We
4COX68KALQ65N3qbvQ+RKkvrpmn5S7A+dzBky2zr2DDG0gxwaGU/lxNpTbyFsjmW
SlKALLvOgJY70w9BD2bMA2wja7D+htkamqOaxtymXbVcj581VFZJUh9G6Q5N6t8d
P56ey7OhGZ6nJ+3RMeK0TSPn11Eqs6Msu1jbkoNt6NhKtCQNsrewz/5rrEWGVNNi
oxUIAeVH4QbrVgW6wxyFpDCJiz1RTk+sFwPAJ5hUJDGxoIN48oEhg3c+DcSJJL19
i1b2Edu3h7wDojBwSkOdALzda9IY6AYSQa8F6k6NkBz8ycdFdfqJ2RmK4ztIoVU2
WaPc5xrtQW3DA8yujrbGy7xZQWd78sXpZ6LfNjCPYYfG7GWi3VL8rSwMGqz9F4pw
Isz9snif9d8LMyPr3N17QxJaLo25ZUrF0BVIZCDkR37X/dNQl4vQ/Ok+6zX9Pf3k
Om3BHEvYx1ykZOmZ32P0Zuvi3XRht6eboUIH0r5PH6TmeEs/ps46Pef41gy/F6AV
cpHG9ocqpt88Z3fPix/lckQEpGKwfYx3R2UHuDkQ9y/nLrFv38VPBrwPsLn4geC2
NDNaOWVPsu8sm4udQmraL7lL9TnkyLYA3WkeheK0s4ymnbhWkiWBoqpfmHIMCwE2
iPPp0v+oG7u7LXBXS9P8b1vu0kJrkf6yNsw23c8hMulOzD6R+7Ep6NsEOj1DnUPQ
LD+6vDOaWj3uIVuUBPlWwPVg6lbp3NZlT1vUSXnQEaZp+1PsxO/CPWdRsr2M7uTD
doqMMo+iz2Jg666QvBZ4jPL2/DO8LNTL0H2w9ykFZIWCOCoQZw9qEpR54sRpf/5D
6wywt5O6wcFjmyGpX5rY7TpITmIrVmb3Ty02RQBwqcPPLHp9hF/GFrwVW78thfwZ
s84fG7ibvxaYLS7dMHEEpjLLc9OCmkPdlHkvaIxjKcrOBhBy+8tSR04sKImglNP/
pZhI/mn0TubJhXr5K5Unhnygz81sQb+Gl8rwcVQyVsb8ZJbByapxYo6w7qSnr6/M
sKo3NjyxCtZjMMhCPK5MkNIWt82+sKhi6ee7Xm7f2zX3K83Vt5yKBwizxLxr+YO5
hBralJG4RFfQiNllc5ldiaXPA/7IixuBDF9F+LQpuTi4G6VIX4LiTeHqDH6dGYGn
9/tXA+7H6Mq/sk3TaToY5IlL+VOVcdsexGZnl2cP+a3QjRDYOdGO67GHhFzKMU4a
EuSfRNU+tmKozrGo15LVNe9C+KyJeXuwXkkw5YOvvymJcvU42ldDkKqrDujPYCGS
PBFJ8V2PfKHOF2FzreoWYCj0ZaxpeWPIPFG6n2cCJ4Z+vX2CE/r6x00raUuQDoUY
83s5n7DRUnkEFRuI3LPrcIL8vrbosEs5BZFpyRQNcu1E68D3Zw64QgomOKGvuRcA
0UxfCvW2TF4qMjeZM5lC0oM5jVjy0zi2IqjwVCwb/wqkdY7ypaqOuLWa9AzGJxvE
zmHDEBbdePNEvabkgiQRQPuNwnb8W5eEv6wf8fsXhQDyDUgSjZDhCyOlC/3F794c
urxmiKU/hbvj0oF0AhxDvMDQlSriUO352ZoIK0eLL0HGs2fD+vJjxToLxphCi26q
gvfn+neWsUSZUX54fqeQK6zKOBykXHs4KUWddfatkimDBQiNYmRmmkoJoEN1RDx2
WWElWxaD2xuW4GYWFNcgEo1s9Z3WVojLkR9nivGsBenCBjIwZczNlwKLaYBTlYMf
DioYnVKGoQTVs2EQMiR81ZNzcsRIB+mtLXDplZaxY8RwO6lm/J7iv2gvqqhXhxa5
Kdnn+mRipr7MAtYqhjIBFj7wXlJEul6lh3GWWxGvJPKCbhyIAZiN4F+bbb7UDJhB
dW55xmJIcIpZgUdmFMs6Yi2TJSXXBFH/DcRhlFQeeaAvdkfUQGS6xDSxpOL3u39o
Z0ajEbjza6EG4Ix8jyC+X6/k9iFp1HWr5wKcPwOFfFl/1OGdBcj8WfUKbwmot3PZ
sMBr0FXG2F1lz1J2CBMZLR/CwqRMwW3f3DYhUmO6pqvseKSEXC/F+N3xBBgskMAJ
WIGQGst+r2T8s9jaCPxKuU45ZLulbwykf7qwOnC5HDCqClhjM6RcSpsBzd6zA74j
segqmvlng4YBGPv72KxoBvw2cACVNBc7uaGfhogLuJ5tS8Smq942QA07Q3+yvsXD
7jNoAPxSdFMvaRfv9BS6hYCU/RdqU8k1Tp/mPst3vSmT81paCbAnxVDr1+GvtW3p
fs3VA0nKhnRkrsmZEZRZd/XWtM15PyJNIjzzAzVXWV/8Q1PaS/uzH/uvlRgjrOBZ
a5wlYlcb2B90DC96m5nGQeyWLzxuBmJeSkljV9ZTf6kafzkZJ93mfxnMu9wxfs5Z
bjeir6rBNi7d0WDc1JVIBkoCZHaLn+CK+zGI3/gFHjZJd7oQ/Omqf+6AeKu3fNnt
2IogycDM7DGj2fL/1rC/d88l/ZeTvWOFEZYZOBDLOIWC9cfOXy6SnW3QBn0BXqSt
fs4amdUB68vYxmuggLwOG8/wWBq04EBX/PTq3nE8IW1RzZhn4mKLhWLU+Ik4f50Y
T2iVYfTtK8cF5/t7CmDtTV3gcxoy95lCxBqflTK97w/wiXs1ev8xTbbg+74jQc3T
9ut/OhOCdLyIPA1swM6azzrU1A5cqmq6PlX9mUfL4DJ7sRn0GlqosGlaDUQGbEpE
qyNck9KoUpGd43mK//HURjjHiGgFK/Nr9NXTRMPv9UjlsC575dhhuOmw/AswstA9
k8CMuEVusKv30yX1b9hBPHYEUUN4JVNd6fLHodSd/Y5pouobHA7p9aCAIBvwdt/5
GfPHaHTBap8UDurU3sB/PIiWMJugaLhrYgQmpgLJqKnTPVmozR1bk0eQ2lGvbQE7
MQlaBLQT+UDUWbtNvl800pl1uLt0mUQTohIZPdkO1//CwHOz4nQYFen5wj2yjQ1w
uJKq7gf6XT+3NyP+eHNXUxZ3dmhbCFovqfmQeyPb5pgYjFOirtnvBoPbJo9AWHpu
Uv/GgrkvERAuPBH4tuCPTPHela1ZovcD6GVaem0I3nBVKGLXS9Vey8WySeFSEbwf
f5dwGquUHjMbgJ+3OfqyximR9WQ8Sruvy8nAY89f/qvtcHVWedVmrL4I2Hm5vy1n
JCGdN9PmlK+/kbyHoQVQ323BXcCK+S4qjB8oeh7BqeqjLQHwLfDwnv4p/ryCVXR9
mE8AUex/D0QxBAqLPuv1QSsPv94Q3JLFBMkncuQFp6woTLGYbwnC55u4xcJNa1aH
sI9rkeY63jCXymwGBdMuTfiatdeAQ2xPLKN79j/yKGVpKs4aQzRmZJOgf1O7lVBa
HvVweeb5TFa8u8F5x7GuNPzvyUouraUR3Eb3prCOYwwQOn+a3r14qiVMGSB18jii
y1zBj5M+wwFhoANas+96shhTZZEzuiHxG3wpk81DCoiQgb+XYq0Uk7jGRRiiTbLA
Z0empFvFYt5HiUzP0phYqNZjmDUp36jDRNGb3IGaSemBaXxIFcE4TY65E05AnPLD
pFmwCMTfA/SwCrJGCRg1QrGUuZfp7meDoQ1XlxRHsYsXn/NnwOBa48UtUyGFiXaa
UxnqBk8qvhjdzOMmDbMutkygr13kpaD2TiSxrp2I5++MivBRr6VoGCaLmbbCOnJb
pPnwcTxGeCbuimhN2A+vaNN9KPpKzhrWer82nbFNiMoUWF7kl20lclH2YqapJOc7
klY1aiOnIRRcSILvbR1DZymvAJKPXjklWR2ab9OO7szjLmMDXkx5nDEmFr8Ufna7
dZqQHPAbr8kxGQoNeJYDhQ7ugc6o6gn3HW4w9X/7VkdUZbEnED0GU0G4kat/kfrc
kcYjUYE0jjFEev9vlDfhQMF+DX4sInkb/YnsLzOBp6KL3jOVZLhmVt3t9KXyvWo+
5fhZjr/jESCHrYdZwwwj0ofLOBY4L/G+44UTmSU4SDLYb9vQvWBRz3S3lwDlqrvp
9ziqJrldiqgl7kjc6l9FASNvoVWAhzLbTT7BXfKI3A3AkiHd8P6NEPYNHLHopUCh
YAPw1Def7L1KRaa7i/mVLwlvtMOhMg34tppAQsvmSYW2sAnSvYLHXmeKzI46YZ38
/u2A6cGQvC9V7rON3+iPkqQ/HRAvBt58lonmJii8r64QgRWAinQIFyuCdOVSToSg
nYlCw9MKjOn/gXcCkL8GFCFRa5Z2cplwlk2rEHZIZ3dj0RTB08OO+xeVNHT84yfh
WR/ctocT1hXW3VBJhIuNs2KDpNShCVI6IQef0ZfT+Rtto65SMxKBDC8QZo0J8wMZ
iBR6FX3PqkdjrQGw9Qy2EM01//o4wZjVDgqkAfAQR2FZgFzyMQHP64P8dhwppCm1
0/Z778zpA68BJ7pyH6+3vrp7dC4i+nGQAHxOWwcV+Xxa5AJY9E4SUVuVOLPWWR0w
iH2gy2a3s8tMwjy6RAX28Wr9Zc/IM3BoE9FAhGehk8RT6P2ntIEX7SFMeMbX++Qx
Rakvk55NSxbKM8jnyY+PYJzc/HgfkNgIs0Q2wJZp+bqWpu9WIZNj7VL3f6iLTZoG
MxTXvvCWOORk2UoY4VpEt0Ibcyme49zdZud3aKnhL9Q87tX3BBG0tudeFrdO6bcV
h4yLlKfm0Qzi6+aSXmemAXVuib6tW/dimHCcBkXT5iDO01m/cDoUodlLYpS8tFIu
CsjcSuxVvBifDDQiRWnhgJqQMwlsuubrqV9YoYvzABtUBtG3Fz1Uss8gwphTlXYx
7QUhGbAqtnA2PW88vlEnAxqgSnwPJPDSFsAKeNG7a7dVXFUjEq4aITgRDMcqVlzE
oQ6oc2mAn0ABBIGQOUtdSV87UYiORyXBnJ6d+zvwZ1mPIb9sK6JDN2ZcIUiFMnR5
3KK9edpQ8/zLv/WP922i4/4QZ+ZY9WX9CPTcR9sBlpV77LHI8U2RXszryjBphkSA
hQ2vUMeqWl7GTrfVCdtQU5qXIc/Lyx6tE4Qs8hgyVItFQ8OjWs1h3mnaBp0R6N2i
g35AyP/B78nqymfPDeMemoSvJ+IzISncHILXVvET1skjXOetW6eNwgyMD1EPMkQR
rDn7aUiqe6ha+q8a8oktRWHKoNpDbGEGIHynfwstpGfUq0mb0WkffaVaVHLleo91
pTwLsO0CJv7VMG/3CdydxnVw1UbutMN6etKyslvUxI0AD93paZp71jHjsJen0XGg
bQNKmJFmfKIV4IlVEy0AD2/aW4O0gJLJugMRxJzJi17BPXe9RX6pOdxK+7CRuyqK
ctvpOdqA7VGv0y29yUwpnpS9jFJXdSnOIAAbcJyE+ZUmpOxr8aKAqF6avJDAvkIi
ZrU4dnYlqtyvFBMJV4zopco+WYRuc674dSQcIDs9L5i8YNElTA4xb2LnRonD4NqZ
6J0Fn5Bgi2vHC79Huxz4/4JNBh1JRmVCSCCcmgeXKvpSkuQasngUZK+XLDIaENyE
02qXWVVkXhu5Re5olrfE89ZBWjlSwzAbTV6I2UGKMthVpWlVHANE+rjGEjPBWcjo
6NB68rRpwBpEKYz2DzfOhwBPiH0kRELoVJxare8R1cPSU8mxQHVZeCs9bGQikQDv
BKxW9Of4Nqp3E1huUxg7CFcgHOZ+0LHOJCe3oNRV+RSUjawXkMwypo9IK/ShpaeE
8i48QllBeSpC49eWX8PT7U2YDFFEaJ6jdPwev36aLlu7Ps8/518QPP53EiCO1dH5
fH9bkFhJOblpSk1QimxLSHB8oj4H9hdh53hp/zFQYju/3YOO61L30KkSbCCRMd4M
qcT980ZyjdzYZH4T0iD1cKwUtXdEmMHkW0XEZb1qdmutdGpo7zOuLzHFZlPURR4b
0UNg4OlMQVQ6WIWnmJiwMr2ejsITYvv0oi8/IlmL2kI8nX5ICdDC1bEXDuejg35w
djAGF1fPqHtCVIgZJ0hjbwn70nLkxn+KnPCdV8/vRWHINqyVeAIFdoALbGhpocq4
M7r7pjg/69lvhiGb+xQKHU5TVfBzWjRQ55ztGheg5Ru7r9RjvGxaBFu0u9QjFJ8Q
gp8zBiymXfN2GTmKTHJHjbjRuVGHEF0QrGEVHhwEEdqv4+7qbLUedOLYy3qKWKw9
8Ao/0R2gHZe61CnFsgby8VWBvPDBNYsjHg96NH0BeST8kFTZ0MNtmPSVRoetzAqa
3kGEcVLRvtP8rVg+wjF7YhO2YAAITTEso2vP6eOyaB+i36YcK0KVC4yKlD9Opg6H
BIN7PcFRSk/9m43m5s8ZZ/y9z7p1daYty1U6rSRdPJxOvb+k10GMms/QW9dfnfRS
ELW0JChM42YyKAyzwvZriiSSEOhgBkxwmSgYYJ4xEmBB7AVUneS1sZakRH319aa/
MLOfhw08dVxAyhlW6JeJeR99hocnQPcfFOnuMmHRlVxGFPjpZQlkXOiHXryC3yDy
BuTxjoYOflWPpVS8UTw8e/uwrjSq0TFXzt3nYC0iputOP2DScna+0OiKSWgJpkI0
R/5fOqWrU55jk+dQK4+fa5McZbfTQkDNnpfIcxucwHM9vU4z1SgDjUG4HxporUrW
HiCw6zOFyKK04v/4PX76FCkZ3xp6aoxXtheaLd/OZAu48WjAq6l8f8aKsBiwcMF6
XLsWbKMW0rnB7qt9T4rdIc0tpOeR8x9zYlmUXsngQgXGijZLlZY6hku+RPMt4XML
+t5IJchpjWSM16t2GVyVQi/jxV2zKiSbT3FTIMjfC6d7JX8Iciuz6b1in7GU3yN/
+2FAjWMW88QuCEpAsx2zqe6gDbFNBJgXg0P39UPhiNUCar10mExGmvZ8zm6na/Dm
ZH9AvpCWxv8yCShs0WjZjLj8r5lQfJCgkPVjUB2kb0DVtNoLTQ0wOoMoVZNGT9Y4
y3BVKigyJuE96fGjHXXli1mZwYXRxV7MJ3qtVmElIdO+56kTUBwO6TH/pP30iUhx
4uG3v6DA6EYyp8r2NDlKzJI3ZHcVHFOiY3pCxYKG5+uaoSPMIUYlv50o4/oF9/hc
ZbFys9jYodGa1z9lsscUH9XEotzfKpt6Dy22kMs6l+5xB5cczkr3J4xqNAxKmoF7
8k0tLDkjSoMxExeD2HBM+5NUu12f8u4zi5N99exZKRR0dJ6JbR/gqDwXzpUv/RNo
zrQH4iCQPZRVl3Azkf6Gas8gq62Gja/FxkT8/u7Wb2yaJr6SoftZCKmcXb0RdCNg
piGw5l3/9JlGlt8Y+1wWJzXzNSFvaG2PxawQ7u9XzHfJMxH9LO/L0N8Wr9YUBjZc
6hFFxnBXKv/oYv4ebbVgGQi+NKgH3ymwmAwc3ltIMaNOdR61A27IfCO/jkkQbgVn
gv4RC2OwCE04Zf0OBF+4+BUjvSOPfGyqIGEVnNfPbNfTmHwUTDF1ui0dUqlnJJvV
5XDV/YffQQaJBWhmwWkCOfCOohNjzmMEgQ2mOi+MVctHhnz02J2t1w2aJB/LXjNf
M+4fAJXr6rS5cuR9Q+clr4LEvpuXsgTkCNJCRiB8oQMmgwWqk7Vse3IqYEsqRa5b
c7Vr0EoZ1K1sST2We/IStoJGexLQShjjWXlEPDAlrZOGvmvk4jWpbvQAlc6DKSgD
S4o3NxAuHrtYoRL5i5/4xF/jN27fzi5+gaelRJoh9wIOsS//YfSCvR2v9agLkiTF
D3hhab3/8XyMFOrz3GC3l+uqOFxk4kidbzN29fd/AbWovEWAOUu1ViMJ74tAiAP4
sNcheS9HUEHqjPk7ZFWKqHdsjRssJY06fMaVQGfHdVjF5YDRkRktU2iS2PYXNot/
QxSwi0jCPtdYmWm/2Srl0WdR5oSlIIPVTs1ILleBmE+3hO6Uh7sgJICT43HHcCf2
X6RJ1fbKAJtePBRcOEd6rh5w3xPTIdv7Myq3HyoHsitb9+E43qnwCUzlcOwhf4LD
cNAsm7jET0q2VhJB22Rho60rvRbiURw3z/1XlP8Drc25nwZIADuUpKZ0C6840GRr
XvoeGUB1Jj9tSh54U6r+KIbCcJ/GpzhFxcAwLQiTqb3R+v10IWXQtnOuX1WcnptE
4zN/8m50VinoeTrcnulrszneABCAM+9Zeb2OeNF+a0x/N4GCDnUgW/LrN2usiK5i
WXpOt5OD0CK4Pr+liNKxEuEm07EoIpesqszLWDhx/IegJiKKtjg9GJLCeYDy9EfW
pz2WjPW5tttV2GI86+0bH+UjNQtM+iHB//uzuJzVOIbbA9ej1NYyDINvv8jzy4d8
KUfyHRMbpQ9x6H3uyiTDRqUA73U4tTWuoBKrJG2To7EPBzUwpe1H1Z33bLrj1dNw
LFlxmZXG0NFjJh09VdaaDxCoegEvvtFQ+oZGJQKdaJag8samNIfgfmDgvGWCE31k
YRFZf3qCTcFgkxxo2TC7tnFntK0CXwoCc/cRFcZ8WqG6/Y6m4+PT1n/jUONXSNC4
4ZdO072HJBC44VZkg82cW2F9RDq20dHUQKyc+zhC/a7aP2MR/HIQ/wTNKZzk+O0u
MqLY0MRxSb6FWkHcQ7RNa65nQDIEh/qnwnn7Vd2/+6ZC9miF6vdqU+Feox1Z+CVi
6U5ZQTnw0WxY1WC4yZ9+GQWexNhui9iPSSmL0PpVKc8JiGGCxso8My4uM5w7jg9Z
sQiIvxc+HAgnO1U/ho+6pVwFK818OYy6Iyd0Js9EG+OoyA8wWqwqajUhF+MVYqoe
bxGSoDx2leyDLjzGHULQPpuORHTiRBRMFrFu+F+YRonOVWzcl9QtMYCYg2ezhYfK
Vg9qMswjmCe6ynBAIHPpKNS/hC/k97HYUT5eVkNwRISV50wCDuc0zmM9TKRH5qDK
o2f18uKqRRzlOZReT/Dyq831V2RuP2bEKWVxByDxVIIrEMDapx7SQ+LqSV07qPTs
aUjzy27HY7CKOdEqNsjwpnKKSLVIxqBKp4O4zTWpXXNjM0gZzMyv647QfiyJTOyr
TqXZ3SqJxu2mnbAXrndOSH8xttFBlrWc1NCdpQvd+vta/WJF4kDaivWQs/qh9cH1
/YqApommtRsw4uzBFbWmdBvMqs5qX/6J3tV6WXfmEg34/BeQiOCmaWtZ4z5itEU+
85MtjnN/G6aCDHqAv3v5yyMyRnkRe4fC/d4et48WH6wYXC78gWqVPVCP3K4QwARl
JmgMPL2+9vKQS6OI27iooG3iLgZTnlWUMhE4qF48G5u0jtpPSPzmOvXXEzRO1vC9
mYUhhBT34AC3yG9zwXe7eY28TFFigEwB75U3hV2xnQqGvZxGJjz0goHQi6AsEPdT
WB5RJiPpk2UhY26p6a3dJmzJqj5/NKdDHYAvG/AxxEjybMlVZoydEkK+uuZvjMvI
a7CCGTmthzRIADPzzpEBMqRlDs3+YauXvaS7LXU1W/e4Z5kWXWtD0FlM7phssu0S
IANKxLwQuAUP7ALZO32ogkwNulym6bMGlzNyOrTO+y0aVAtDuYyl3ScjQjiw6ajV
+N570p0Sej/4Ltzcb3ES+UUXBO+m84BqC2xME+2mvTGNiv255uVfrayMqppcKbC7
zyIrznL+i5ILkux52UVkzvouK/Y99Ca8f251BcZ5Cie0BhsDdg941NaPirr6zcH0
/4Wv2Gopr8piZ8C/aqPvSdEig2rqHIepXghRl92jCsYq8qlKs34GMnr8kmgBmmvW
O14fW8rgxB+CrENQc/iykKvHSSTc+vx+PME1RiUko4UHQZ9qFLioOmEm7nOwowpM
lZEzwCQmrm0fUk5xJBKNla1k0cvPp47fWiNT7ERD11x9RlOOz1jMsCeSfRNXMZ3i
wgtT7nw+TJq5GZRc1zwjNuHoBXTkBCW1UCYJy0PoVvCMQD7+82vq3UV/eWKLY6BY
iB6r1pK9apdGKMub8m6unodTF2DPMD2C/+nlgR/z7DPZrgi5GjY0xmpn329vt12o
1E35hZo22svWFrLmEOUUzNiZ7xC1gzT8fef3sCLDStz94fmNXCj3F4u6867v75A4
kVbpVME5elDm/NlnucXSFN5U8Si3Alk25xYCBFGPUJuXOVI3xvuLRHrBZxa09L91
lOsFmChH27d5bsyfV2dnz/pN+WqoOzByR0FC0et71WICsnnMbwXS81p/PHjUNv26
TWr2WJiNDK/fHnc17gH6k852iVLz+cv2jLnwGQxvc/3pyT4YyCj7GsrjDvIHeyDJ
ye5XYZDLmaANMlV2WbI+t0hHiqOEzfz3mZpPHDGlTdcvxC/4YJowfDW0ibsD/RmV
lF7+8ahDkizCeKRFzAUsZ/DSxxtXoS5uRHG2EgWCZBnucIZHeRjgOTaLUBoKRMUw
xk0KOP46Qo+231UssZVMBKou84eux4pzCUF0UGSLHvqxbBvB+Fl1hdr7/kFlo547
h8CQsMn5k1gOd9BRklYBVwrOMNx+DS9Lbn+uT5N9h3lFnd5+4SxQyBISxgayTq0I
CJFuYM+4uEjQ6R8d3DCCg5MXugJz0f5jpD3om975I0PJouepb369/BststhlmvAO
eA6238AtMPjkqeKEPRYpVLygm9meCy2vSKCqsmeYt6HiJQUm+WJM6wqI8zU8uPOH
9ezogCTa68WiSxv/Aby8NGTRzXmCfrhMI1nkSA0Rkbxata6d2LnzaT8BwtmS0pBU
hpQ6seehuA+paSsIMFZL2algVAoI6WpqJAIIOve+o2o9QcZj4dpjSOu4BATM1gBo
bAlrB6a7o+4tQTsXiE2hvV7yG1TYFFSN5ptCL/mEYRj91hBAsM7oj7fC7TV5N8In
o2Mq/2Cb6Zps/5uZZvIhV1yHCqUdzg6RgKa7KJESCLQTPifaIYM8Udk9jGz1JMJI
Q/5Onflkr/DFUZcnGKq53cmg9S6HL/BxjGZO1BZ6+3P0PArFIOzDChE+yqpBHMES
SeLPSa/AXG2wn4qYJL+D5mfMFHtpiaGkRf+nAwV5ZEuw2ozM2y7qMmyhf2oaIDCq
Spk8GYOlU6XuNxNeiEj4GuqDHBdARTH2Z0opAFt5tUYsS8uUpI5kJ/WVwoAV4woy
QBLXBds5kvVWpdqoC4FWIchmbp8NX65OUjMNcg9jvzOqqOrjjLPKvX3nJt517fPr
YtVZKAftjtwDglsnDRQXgSrtp+zyuXIoRSK8Q6MV/6KF2cD4LBg24qzSs7ppMXn4
cGbHem76ZaR1YXUlHmvA1OYUqGYUitDoralJSySlqTUkbNcyhj9rIokNyJE5g3LP
8FSBpLzo0XesVyP3QDUMLRZh/23RCjL+b1eKxbk2OlcIMxHfcFD+7j/LG2XjLRcz
O1qt15+ACeVhSnS+UJ4s+lrlRpFojzQUFgLxDk+vMu7yE2lm1i4KW9nqt9XCwLD8
J0RaZ0yzATr2MccoXBqQ0LwgOjl1b+7M2JYSkY2Qb/ClqzS9z1KvgEftJu7S9lMq
qKjpHwUqfzhplYO5FnsNcVcVq8/6xc62CyMUe9CnDb0tPdr1zqIeHuiIe1HCFbPt
nqdWGzS6A7PUcfWbrVLNJGkovOZZmPBVx8jyKty5GkqS/9twUdOOPXflPCQ8FMRP
+zL4bnwavKpI+OFRpe8vIUPtt/ldgC3wF0rAyjbEoXpK8XRyeaOJ3Rh3LCYE4bgW
hubKDdQnSnmKUG37kkWIrvTg7fb5LfqZNj70/z9r9mYOKl7gfJupIhZEeWCHtQ7v
sLTeR2f6xXu92SP6N34lWHWFq7i56C5K1ioXk6gxasw07w/a14WayTKb840Xq1U2
+rQbIWdGhjb3ebSZrsvUhXMtHQW98MA/j4TXucWUYkqRjLNzLIfbFKDB3Bz58xKf
vTid7CB3RPpO8CkpoFNzOtLchzEaEavdG5YMEQMKMtEeKKy/4cTW2XUmeBeu5sQa
Ixalhs0/3WFIRcTnB5fwZ7V5Ia4Fd8jeMQnxRMIfWvwYbQVMSRCV3f04R/LE1UiH
3QDC+qXI+Kh/O4K/KCqdns4d3SRyxffNzT2DiWZuPsN5gRZi/4fovsEt0tHNb2CN
rVk1khNg7ggBeVxdap/4XjNsGeVkkzK8pvNEbfNkvjZQVUl/K2iS4/Cm1dGTGfar
gmBjVKtdWk4Ofsq8JVEIXSMqzKs2KARhiKwk5ry6gTNmIlsjRCXRiBsnphYT/N+V
S67zrJtKaehvKqE9wfG8T0JaBnygO9sTCch5Z0d2X7yfz0rZEFMeYWzYdZyvo8by
qphi/AfGcM14ai4yVAS8keqrmlBIO4AJLomKLWFw4vFvMXLBpMW5KWf6G3KLUi67
qJ7ATRKJBVK4ziNc9k/LjzcH6qrXf8zOQho6amFPshwf1eIN4E3EJXTCG64G6yzU
XOu2jg89lZqbbUQsG/tH69FlpsQyxAdKqT9gmBHVV7g0DfjZ2woPdriWS7qW/H5p
L0LkbwkST7KYYtbrYdMYl+ByzALoF1cyjkkbeVNOlRvDJW0sXSWOJf8oppnGvQkX
wHlT5U/zKRmRrI/Y5vnocBo1znlmru7Q8vCjkc88uMg60XEM2VGXDj1jACEj1gOF
uC9FzyRP45Yr11XJvDUiyz4uYfaS5KCMlDPZ7KnzIa91eN4ayuI4Zc6AV5EDbalI
ufe9jZ4mDGBnu3mIy7c3TCpPBZAhkuSCrh7XtEYRHo2IiZpSYnzdIrEVlHpBX3j9
SOvbHZPtn+usbM5/w3kVY3feUo51TzNrl+NkHrbHbJ1E1n6h8eHs0q4QfJfuRcrE
Q5GwcgMeoNLcAfDDncSdkxyJ1g3GgHLZtHYX+1K2eAvLvNBzb0CCE9SN2XI4t+BI
W66c4UnkO3oeGwDOpABZYoIZXedtnm5ahlNNvmi7pfQ+U5uxPrWT7hL/b5TXKY/V
gWh1QZIyDZTPrgFr3+hkhi5cW9JYWuaCvscM38Tg8zmQfW59X5x12al7jI1b23yX
en4Z8lspiUJLglsvOLNHK94TujH42GNEDM035DyOcjtvI+XqxnnedLlug+2y5AKV
yhTnQT9QKuMMSnRJ9cHCrhbhTHULhHam0E688dIYzyuRpiZDv7A8Leev8g0lWJsV
y0gI0Ql/zXkGQOZ4EoBhNZcbmVJdkoK1owhBeWWlHgWwduNIYHS/YsixU8ABLjbo
0MZ4IP+5aPr27mBokxQYQBbGeNJIheUrZH+qMHMS0VXCd0M/LI/BSiaLMPX+jivN
4HI55ENPKnKQ22kixauIBs/OzJxhGLB70A+1wegH5Ab4j5lDnV2zPMk1KU+rqK/O
nkb/i4BuO6JcbTyEOTGEisfk7m4QLRp5dcA1ZHal2yaPbonJRf+IW36t2NeEskz9
EZ776DRMzOGcPVC9sbAeKSsf83l9N7fWyS5w1/Lqzp8jJl7zZsOygrqmurhehZ53
SD4cftOaf6t9yeCtSqo3CJWzzVps4lKwpYyjvxR5pta1J+FZTUmjJ62oJglhQMFG
rdI7amvsoBcPH50tC53N6yNLpMPcnlTB17w5TMyxxBW1qt2UIlZudeca7pvctrd2
nXbLqZNAO6FMFyPOQouCZUZxNVEH2w3H9Sl7hBNXowz0qj6AityiLfnkJxEHz0sm
7ZVkLxHvaxinuT0YoZShhbUFf1QoxwQOeKvK+agwCG1yR6c3BSw6DuA2k5pVzLUz
erPPfQsHtXKZtStbxCysmCp8rOb3UWA9NLwRWJmYgq/VlUwMmDsJRQb8WnGL+3B2
wg8KG2Va4PhzrV3LdDePqev+yWxzg9DvwKD5Tp5Hxnzb8c+KnzDDEaraVon+6x10
QMeSd4Bgt1OSljat3TjyBqAR7IrnP5IkI0P8pDFVdRyO0RhjKMm7e67w144teIql
jg470csxgVNJ9AUKN4r+aGS6vncFpQbXb5C5WuHJLaQIzn19SXdVL6OGyaG1lPTk
ZcLA9eE6sw9XrbqCgQa9ZFZ0UYTl5Di6u2FG9A16zB5AnuthaNhQF89pJ6GMgAvY
ZN18nDSccAFnasEZNF/A3JWuAKvTroJ5srsNaEjC/TjPSXBrtSSGkCMez0zf7Z9z
DsMcG+ADTdTqyRIeSiHBwbZwfDrvcWRdu4/y8xJCd2X6b2CE/D9p91sWlMnuxyW8
TbnFU6W6tdF+6SCTYNGPUZvgEyYyph3PA4+ZnDqUNRwMMytDukyiSTnqZz9hv3v0
jYmt5wyFMd75KxOj2bZ5zkUFsz2Z04soAihxhfCb5QNn5Uu1ih2UbwU1PxtbpvL4
xotE3FT9SKReUVoeKI/ImL0u6I+oMZsYKSxLJG0eqG7PZt9+jQ33J6kxi+WaJRCB
+jcXMujWOsScMS0YEiTxUpTR6MA3Ii7tNPJK4kdAwWuhvmuhnKnI28+FRbmCKhWo
2pCpeO9Sta6oQoHxtVxJibpUc5NkqsYwROhMqz4LFC9d+aiZiY0cZX7TRrHlfj6E
psk/3hwiVHEjU0ClM6VIkIkHN6/6QAKOMjteo6jp+/k4/owcRY46KeMyl6CleRpU
e8cI+6UEbnK9qWU6AEzmTPDk7GJft/OtSd5KpbzG/GCVmCIp0GewG+AerSJ+mpIe
0HGUG+XU271BYQJ+FUD4zgg4w6MOCQETGTZE3paeR98jQv7wV4+F2kpU7qPy2Hoc
y7ae7rnKvR8u9KrgxKO7I7OiFKSWgObfDXLZ/W9eoZgw3FxTvK9NiD+y0MEwuePT
oXFT6368m74JlhSstaZyGBFmGt/xsrufmLJJuiCuRSifZtS61a+9ul6bFn7bPCym
xApLegcbfZomRBoq1P1C4MCcKqtqklgPc3p7hbkIZzCdVh3tORmh5W5ffYczx58I
c4ZE1P+k0fcchxRMK0xnZkCnMRPYS3Fd2gM4fT3TpUhLqtBJqUr5RkLp+eFwemD1
7OWp6hsblFds0zs/pHH1C0nGDWbjROFWHbIhYKO2zUmd/0L9bbs5mExyRqsparqh
du4OPPMMLZnproNV+icidHgF4oIAlfWDJdGJEza7vxnit5MhhVFzbq2JTpACVbqE
XyvWXg3a3ot5d2tLMnhiNDan4+f+oZ8o8CX1yygRXg8U20FR4u9mHSmDOpCNIWeq
aiG5dy/tD4UqDxu9+zHRBfd+DFPTE4Hu1zm7d6wluwUCe9wWZoxpc7Wg6g4CEt4E
sG3Ztxm2nMCzfPth3ea/su89jJuuNrAE5gQJlO+dxmE8XGfx61hMT2Au/oJxgncl
lj2K/4kXHiLLi5t7S9g3ezNcRGuNO09nX4ICI3l3cmsb9Tco1IX/5mcep4LiMonK
fDfYfNoZ/3Ctz7xakh5iNIrdD4lsdwP0yYwEgJIETM5fDIq6WxlmdxeTvryNHnUI
Pe+4kjr+mrl0VzogRvGcdW0pqCt/GA/w7QJLr1IQi8Kt2UEB8r5oNRk6Ne9uyseb
kym565z+h9N7fkkuyk8cGUH5TMu1L5M+heGnpRpPud5wReMNyv1bNPvKmlJi0WCz
bQaZQRECQBZoi4FH8A8bOi5CkhAWFK35pYoylcX2wXFQ87/vHIAskiyq1BHFr5q4
7Kz5lV+L2yDtjlg5502UKmcuF4OOdiDIULUQsEiqSQD9hbi2HI0HRsr4R7Dxx8cP
vO7qebLk9APKsI5qoPOpnlhJHoDD9nlxTMZPjaaZhPTuRGCIs+OsoGNsae4DYrDL
F2ThD7AvRKVnz7kXbuh4qUC4ACREKQGghncu6zyd5qB3zzmSP8HeSmZEKo/KvQNi
OCOK5mrUkazfM+hHQYMV04BeX07qgxPtjxbevNY00kLiHif8UrmM3RA5DoctDKIN
lwTAXevv9lw3jEUM9cV4bndbDDa929wy02sj8BlMK3HLOALeQb3gdSV4JIIIZQ5h
UUI5xFDSQN0iW6SKSwS9FI+qZYP9oApyvpbz8tWnGcaA16ZZ/ddgkXwBA9dJ1GF7
QzFiGEAgdmD82AzQRQGOkop7O/2ztP7AP8KSzSu4tP9MPXm1oGxmT+hrBI6DVWHU
p2pJlAwce9CD365VKaeFf2621ljDU2Mgj8qTIbLGXqIjdS1ynz8uz9IePZ6nIGbK
+zhO82k0pNNLxiRD5YRIlDQkiONphl4vKnmbbX1HBGQmngMOC7LU/n2iBtBFIlLQ
zox+yxtjzibr8HvE4hfMFY0mGUpcqJ/u0Xbx4QHQv5dz0gEg0WTy/MctYF63wB/z
5h5snZ44I+hiIXCpJuFZl802sTCGRCumvrlbjeccCetvB6ARXGa+Q2HccvIclUYv
cO09NqavK898/VbRX20+vHEcSjXwIs2oHv2bXcPoMjdlqYb0ogTjIR+8BMrheYER
Zzewu7GGN8fArcxpzN+g5M14XmlcblWmc+5PuYjq/EVW3nmKRiXgRUwW0NnyAdeC
tzQ3kHfISi8IpFeg4f1OspuaoBopETVnqcMKzXWcq1ui35MCat+rhYZIB/Dt2a+J
aBinwqs/kd+2mSEApc4fI7kPAe5cYwvp5rjCi8AfhJLfywRNUVDvK5cFJiA5X4SB
9mcsuZka3wZsj7Xa/PN6QySMXljt81x/oqgPcajIno7fusU3TM14GUuAOERe5KGW
t3nMgbcQVM3Pijhyp53Gs19MKb60dXVN+PT2TJIgJ/uwMUUU1YkuR7HhAtcWzb+e
KCMQGththDsc9RNBRSrLC0izFJ83Jw3WDDYVNlNR6tHM9a1e6QE2nbVA7KSXCw3t
d7yZqJ73YE4jh/R3AnB6xm9kCeNuJDiQkHbqgl4vZLwItieLjij8aw+XAxRoc00f
C/Rzi9U7P1mPUoLPtyyHeus0XTlgx70p3gOeuo/2rI7Pwc37lHnMvtqNGAO2EbQ6
60sNOXyka7B89y0bpx694zWIU5HmeiQ+3KveDuBaAlkCwRaLxVJYfCqsyS/mn7hC
rE89KZxD4Pg0Y4UGTf5AZZn3LNMY7HeA1VsXh1dvbISTT+h6fZdbu2xDALmqsBti
ZbdiX2r3XBzSJ1ffFkLnOcWaNnERtSJV8aqa6owwFY2lQSKQTfmYA5FnteANhf8m
wR7xO3H7yoe+tNP9ab6CvjqWcgp654IXZP1jg2b81X/1tJuk61dx5/5Vh00Ky91i
dbGX7RdzrliDkvTEZ6rs4zG2ioWVgZ2K941jmd8vfYnAZU+gEY4VHzQf7+pbbnkb
tE+AqDWefYrLxPLBgnNJJ2WmQuICKENZ0TvmONn2pc353nefJCrSiYRzfSq6guSu
wBa3RWqQ/R/AKODvd0SC2ug7AXDSF++ZisSsFywIN1iVeTOn4nOW4EUoyiyLjIst
iM7abRVh+l/WHehWP+eP/Y0dM6eHvzt9+XHz8SEhvt2ZuVN8gQABbp2lcTKZHWCn
i7B91aNJO+A1cyrViz9IsLS7VHRkCOtZM1FavZvPBbjWapMtJxAQm3JRgcW5mSMo
E3wZ+65g8ICBUIzpa36DOQreLiDcaDusTp0yFaz/AgnQ4oy20Blb0xIWnrTFAQOA
DHdWLq4Ou8bYFnviGH8zsAMIujJSsCv0rXz1u1Mj5Ci7efNaJI8ODiUk46stOM+3
K9kp3NX+xEZNc5ZOjHPISd9+ut+DKHt4jbMRWzkY2+JFjt8PubmRNeoEWz2OqRUN
2ZUZJhV4X89XkRMlfnDXLT7JTMzMSysvi+xNgaCLaqAjDyhpSF5z/1Mnvtb/g+hX
/wiJqWIttidMkv6XiUgYg04Ug5u9q/kOgwG3duWb6MeN8qlbFJQJwWzws+59/23Q
Olv3W4zfqDWyVNgn4CXR2lwQ6sjOW+W66mggEztTOlwHDNhnk+7eTVZEBGao8gAf
37t6jvj2zRr/oQBwzQ53mRYrG+hQNPCnjFODmGGOFGn3GdAhB45qcPlZs6itk1PR
IBIbe2kaZ0yjdqtpkwpML+B8YAOx4HlibLqspnPvnY9H2VcFDnUL72YO90S5QH1U
ZLlBlWsgqg1KAEPoZ8zvDCaJDCUTAvBk+Dm9/hwe3c9HsnqnpuUl2xlVLZpKwZqb
AoSETeOUk39oJMQtE1/Bfhy24q9XB0tcKCPAlfev2ngoPkvi1qUnCl6pfGbgK82d
Mk9F/jSMAvf46EK1HYwjKxUloDHHGMnc9Aq8lFJCj9zQ6S+/UQopPGb7hGy8qZp9
KRDhte9kNODoGLFjgR2utQfupfqtWTa0jUq3okjQpcyrnl2Py+lS0MDFKdP7AMVX
jkhUkJMEicRdA/+g2nLp6SE2TDEIQHqJM40UV+lEXYdgLy3j1lJl6vU+TtMs7vN/
GWMSQWlh3m0n78e9wS7VdIUPa9XQ4MWLk05roblbjQfiCaYp8wdA0CUjMVWxYL2p
3SLTpzeu5bz8JXNVDYQLCQCpk09e4h3WG33VLoMEvZkU1qNwyWFp9GfTs9p03kKo
wEF1BcUSSREMoXJmmBFvalRCkBxNtYJt2RW+rDP5T1N5fhGRyeVNrGYAIyo/lA64
bATciRfCoVNDcaWpJfByMmhK2HDt0/RHEuD3rFmQItDhvYf9DcDXWqOokh9PssTp
EVX6nKUdadZ9y6XjvrQLlMsS6wM5y0N5xgC7+AOpFsNChvjyv9i6fAcYRxSIkgu8
EwoxM83JuQQpgbUuGJhbnQKYk4iIbGnEH00XuB+R2DglesjbsoU9dO/J0TGzFp9y
hqB/lcNhaljcH349kxywpjwHY28JfdUZ1aHBjU4R6qu/PhLxnCfqsb7h6yMBoNWc
O7YZtH3bIG7elRaBi3VCBejeN/qNathRBVBJenL0eY3ppKnFwX6pqRuaU9kdNDcy
TdGsOhwO2RssMhJPfU0MpUBgumEw6oZ/3YQh7NpVizWQNTlxtmfHF2HvrEF5tPx4
7EeLqB7EDfJsszT/p+sz4lZNmj6Eb4Furovg0RNcEdxfnmZtbY3HeWSIE3ZxgQBJ
ViFHCxvQ5HrRsjnc1j9a4ygCSdS11Fx7DXCkcgJL9L92i3p/mZnJDdJtq5zGv3bA
DrgqyxH/bhXYuvJkFSRjQXwROFQgs9NMdFWb/zdUB+p4dO+pCN+V3vanNXTajd1s
MunmvKIcCiu7GOkiSwGR56HASnzRbFlB5qNLVOssgmJd0o0k2NyYqa7kJZaVbLUL
lVp8sY8+TKPZbcwvKv7jnoh/rgMft7s2UVXL6MyK2mresq/YNEIiUCWf/lRYb/hs
NyvWuNf077Dg9B6Fg3HhV449l+1JxFkZbXsePSb5wjshKSr8eiw9X1i2Pk5O7yay
w7Nl756rnk1kohvf2rXWZ4y4yvx3VqVm/F6AtDN6bvw0zsp159dxvGYGtrPxIqV+
BCXMZ2/hcnZz5wiUndT8GmWtQRtr6h6tt5bLmFT8RCryDj2qCubd1uesszr4VGrq
QvRv6DHSL5UJAjqtzMy73GE8kmVIimqI++JjowXBEDzbjm8eAFSUGmVvj0bjVxeX
F0hH6p22fSNV5TH9vcMviResK/kSjR5B2CsDitIV3ghbUN1qoAsYulEJM3CHzYv8
IhFnsZMrSMfNZl/3ajMWD2FaZjBO0oPCLvBdH1ytM6rWgvZczrHXFgTYqG17bb/x
jtdS6/mzLMEBdTtDa/nJmPGNqcmYWNB3/qiea1HfxgVPkWzEqclPzu1e170ckCB2
mPSO2fb8JYn4ed34othyMkeJkfreiNu4iH6f5HOLRdDPO40JGa24DmqfHmQKLHCJ
gqjvoCI6hx+sLk6cKpirz82CW/xVQfXNf9uMSW+BNlVY8KYzFGtJCL9ek6Q1yVcV
DckN+eD5VC0vdSznsF0P5ehftP9SfTb82jFynWEC0QyyU8slhHY/QHM48LtjxJUN
OZ9266TNbtm/vJOjQc/5EKR75oo2PpGeHwvCsib9KoU6I+vJIatSAVxwyPKzAOAq
ULCkOR6WAafR3cj1IHOg2Z0k8yVD8kS4xFJ/BD44DF/bAWPH7Uwaa/0xYUK/WcZl
EtGdKAV/gi2cAzzbJp42QBjKt8VT8tytiLior7KurnjbysDWVNIYGm1JprH1chz3
ZYTAStu+zDkMxFcHa1B1b1wcZAE+Q/ue3nDpSnLGDQsj7N7oNOnjXEWXSkjKIgGE
k9qwxfb9ZkRLpXYi3eaFMC43Gv70pKQsLe4A2v9vp+8BnrsJvGX1u151y/Zj+I13
WBg6lk7QMfQLhNVlSRok/V0rmrbk9suhl0xnDuO1tsVUes4H+TKIrcR2u/aBymnN
uOPZqIJGDfyCP3CYOurR2FcQB/cXKxfQPIYvgsnD+OIzoKneXgyQAB20K/OdEH7U
0eBBAMo9YeMJS1yU4SG9eTO70yedwdE5TU35luPq0bP4MCgEqFuqrh/gcwDq5a5K
ZW4xZ97i0OUTKhjI2EHqsPfBGuzNhryF3fcXWoHWWvO6VK2MmFXpJk/0UiEo+SxX
ZSpJvAEd8XdMWaoc8XJXbOvJDB9puYSlQXPM6Hz4kaL0RFASOjgWScYTLWCc0Qkc
kbLBZJAuYhUIukbzde1aNV4U6NlPzynkOMvGI+bJBi7NlTxieBSst2LmQ7ly+7pf
979ADTqHCU3CNUtzo3RlC3PyqU1eVcuG+JC5kxxWCJrQGhikx42l3ZbTC3UCeGUw
9XMelAJySKEMkPbrSvst1P3hpvbbOHkHhCeNnISMvCxNSFIbRSwAYS9AqF42c8+k
5W6C9TkuhSF2K9wplA8Pb3oYkXAe9t6LRNuf9JBnqHNflobbjC4aqESclwyoWg3v
R8JcHu1AJc9CZcybtkxT+m05/HEX+2lP/wn9cl+sgkFliweM6SSRszS7TPzJXP00
dCQuJNDivH6WS3fxGpoSUUo5pw/zDq2A5X7ddmGATj/OpWsctVSjcJdH2IgK/3R4
WWt8jIjT8advlJWDqXrOL7sAYm0qhi6mNZU+iqNd4qYYLhR4APxcCpZygpbmLYgf
wxEh6EgAHJx2ygkFZbzi8lS9ziFin/eAJpB0dBsehZIJ2+HJfCqP9RP0mrsR+hpQ
fVKxxzkXtVWANS4jTxfIoKsbvRKYjVhjY7x6JprDKaFbdi8LT492HYIzEXFi0m/K
UBMXFbQCge93bsImSl5OyoNQIR0j2nctyrfLH4RMZVf1MZYwEjiObnRyG7NOsKYS
04wERh9pN9rF0UdvvOKflTa7zjCQitQYjKau9QXQC6dR+N14tkWButzMAqp+WD+v
aHaNY2cOnIG1QbiSrH+iLZXwU5p/ZOSuohzqv5iAuasEodrecubF/UJF3UNt20zC
gcg8T0tcP7u3osoxO89iUNW22n4Kn6ZQqrG0uLfALqJS5s0iI/9d859tXoURSIj0
d+ukSarKPU/ItJHpAAkJTnVeuRKiuIst9wkXtZTMRgg9H+2Rg8AIBTU4M63Tfr//
H613HXd8FRO5ktX9HHjaUUuXkWTkHLxgadt35JQmTZbKWX9dDxiRM/3aKQeujWlt
OSe02Ae7nfvogo+A6DFAamAQ64kvSpKVb9c9OXGWw+4DCNup++pu9WEtrXewU613
jLc07wU5GT1GPWU7yI9qo5yFtE6dIoIJQLMvFBKKbZGCLNJkb7xMubCQso3JvjSG
2Bvnr6OX9gPUSxcYGyIXEVS0Gkwf0pfy2No6PGXCC6HOAaavWiFXi8zZgaGkTxHu
ddvUg3l9w9QnUp/taRjCFDynM/hkjnBP/57X9gV6DgGD+e70WXpejuD6t7xSJ6qA
JtX4iq+J+oD7YZxNWkT+/gCSNf/d2F50Ft8VHTDgfKk1rs/LSQU9UC3nuem9IHWt
mXUaV4Q+kqDFbMgY7kQCajqyWhTZH+Necn/HdbvxNkPWNgef+VZr/8Wx8ar6H3Br
E7rLtfsQOYOJLmShIj/phYaHqc42Nr5uQBzwc4Q/toNw+g72cY4OKKuRja6qinU6
3S/kH9r5IFw2UEPHEVGn/AjTSNdkVtxbj1+/2TXnx+U4Okx9Ub3kzBeC9d5bxY+E
rwZU2JHfVPiTRa1ZtcIrMhRvHBiE3/PLsqFUyeFm3WnRSjwv2+eDxoVVC4ONbNOY
naYRYMihPw1/PVCvGJpdx3wnQ4mQvRGGj+q/gNCllJGyMbVQMMoU9/BY+16+55yb
uDNeS4uUkbo5sXpfLAqIhTbvKgUTJ6rnmr3OqkkXuMhQ3JNjjJDT8zHpCiA/zkNn
Mo3F5G478MN11kKsaKH8+7Lv46Ao/lnWWC9luo9zbaMlzhVzQ/G9BjTwAGPhLRzl
gFWuBhvgp5gjBahQ6A+OOgsq76E0xmULJN9/aj4WWXBwqv8JkfyZeSFmMeaSuJqY
Lsr8hONMqGEBBjD0gC6AIy9TZcu1Chs1/u7kiVBkyGSBZ8RoEU1HUy3dld4ZX04s
BsFM8dbzN211GjhF6OIjHDKENNtTLICODEWUghrnVawf6OcYUlxMJ0blq50iZ2Uv
Rb7I1o+diZ8c1MnVKnVPSgKFPwkElfnpZy+S6gwrWWa8n2Mcok+7wcsOywOEs46M
u/xaMQ+VoaorAZCAYZ6tlHtX6TiP98EoIijY+xcOFzlOBAjKJVGfmmqTK7JgdzYJ
oC0EPuchyLqL9dXqYa59r4zky3r+cW80/jwfM0zQNGimvuV7uwTlYGa2WeH1hAK8
78Pyg0i8MPpGcDlcsPcWVRxwJJddF/34EB3L0+iL0IAfqOVK6ndosDlDHqEhpYij
BjbVOKyb6p51pwEKcaDo8/Qu24o9HUiKh1prj8qZhLSvnhswRKLIg9xZ3PdHD3Wa
qiuBIctx7T2N+7/TLZ8So/GGvyk+OG58M+veaBUsJBEMfaP2QDItHW6Vbrdsoa9/
zB3GRJaS9E6pP9qpi3/jSc67TIVjfr6DksbYQcPKGG2leLecpIempbgoBzD0khK/
8MfjiPkpxcFhSml/aVn4JwK4dcWER+brVDnjewWHU+Uew4SFWFi9D0omAFsPrX+k
pVzfg1GLWa09niHlKJgpjpHX9a1r7SQGF4/tMsWop0Vu4/zuwI+YtQUzw9M+iGd8
SkxEbx4oIktE2IjJfd75KfHc8Ckd8K9Kzl6tevcVxzvUwRl8x2iGREyhsM0jUHsl
p48I4fH3h/fJYTgmJCvORVJF2CH3wuxPZ4BB3XMnrYh7XNM3cSaNqzeEamuBkXYu
svDl6GNhG+4s3+qldPKtz/ZCAAopEhfaFy4ZhWV6pMxw97E7+ZqX/62wDN79KrZW
Q4ASpLW0OVS++k2v0ClcZ4qxvHnzVhHs26bD6do0cptoUtF2zrWmB5fMQUQBZaBu
cmik8EinqoutEeXeBxDxtXW4leTzfifo2WYJf0/4mV7PFEYlE4mwGxCuGXGXOJuu
kNP7QWLXvhinpiZ69enpL62TZblBmPtwEpP6B8fx2kIwsCTK8p6OXkzhdtFibpWO
3HZedybJJsUhoJ9yD/zhdO+oOy1eDNwezbHIP/gyIgtcNK8nA9Ma0cqDuH0An+l9
aIRDysRFIB84PXxhFeWi07wkcafsqTH2swXXOPPvp00XwR84Otqt9K9yb+P0R/4e
ZfOE00dDOJjbOE85RUyHpEbDLyk6O4/0nQLpk8L1hCNELjrdtTsjLIdL6lwS9S+d
+6mfTXEJHHb6aV2Z27cI/EmKqq/HtqaOCVbYbcpnk1UYWFrBU6Dd5E+Yny63BIC/
mkjblu6iXwnI4es5gzrQYGIQgkUn8pIDXgjJ0ybD04tBgvqD504SlgPllS0TuPac
H1C6faJsNXpocTt3SDb9X++x9Apj8eRKQMRxqQdw7cI4gudDa7pFVaGrLp+4ruP9
SwfLPdELhZqJ+7feMRvABkj0ssPBvtz+fKkx73PDOL8t0vbXOGlpxD+vicXFmVoD
Wa7KAuYiHaQ4qh5M6BJLCS1ELcGV7OAyAbOEiaMZaDfRtvT40FLb5I4T3qZNlVkG
d+fHeDq/vpShV/0ppikSWu71plaqk+Cy9r5sveyFjsgVI9GydLgIZ7uN2TRFqpCJ
LiMSFMyeplAJCL9xNt4m/57vh3Gg9UkpmQiqQ1a4xDd/DxOD9RZ3ouLybhiWTzqF
Adl8VnUBQ8QJ1fa6F4EwL8m86RnBsmSKIjuxu8lOvFH2iLhVfgslcuMW024SQZNI
kzLO1F3DWHQRCGY+cG+QvRDRt/mYShT49YAZtyRq1o1ng8nSiPpW0o6Jl94WeIN2
8RIBbeayPD7eFdeUJChk/uLv8qezKpNk1TsUMcEhc89KZ0WYSRNg7p5t+gULJ8cm
8DYPAd5mK+Pec/bTMc5QfnNrfdeT5Hk7Ui98E+blAWlwaWdK1w3sYX69N1vp17pz
NVjdPKYSTevvnewhnO1ATnIAauhjU7RAYTuGPWMuy79nnjDXzlmFhChSF6xcvqS/
4Sua/cZQQW6hTv8GeiKvbj4wRpAIeNYkA+fDwUYPxjyhiiwZFs+B2LBaskkgfZZe
p9vODjVaUChpLksTqMJ4wuXcZHBBE3iKM14kaaWhAh8WbQzPCh+HYAqtFsBAd7qz
2FLLHMMB+O01SYvS1Py/JzPydulVCxFzbXBqb0JWVxNx1snSyUAHoK8amUd92VO8
JSapzqOOx4DMe/GUK9SjCUxTwZjhgw/Z9zf+eLpU04orrVxYdp7QRSqXloxSta1b
erkL8Bk5APOh44TTiBLNHJWzczQnfsHWJ+zU+QIYNL42QM2TInP7jBQXo/vViqeT
fTLlb11n+U8dSoDVnbDZU2SzYiKKTNUmHvIeJdVEfWNudJEaIDVrL2PXmSxEqKCL
kkFl2S2Lp7K9cBDYiTlkIStc1S1mqTQzUrf/61YevOtI56aZgAMKZtT3zwAIXDLW
8snHT2ida0LBZwhlUjjSasJoodRf2J17TjOymAMr5sbt2/XLlBDh1S+WRM6uEcYx
KH9XeFRTiImrZx25VmMQDFswKaDKuchCzNV99LcbWbY7EJi3Nil2y4toJkQC72GX
59jI04JSAvrBKS6X5JSVgk5RG7lzYUMcctmWz9D2gp6oigW7KcKzvmh9nCjZZLWo
oz0m2paz7HRfoeYLzAykoBlprPNI31b+//ax8kZwcdLIMpyqtquiivAJOcL5xwvB
t2BfN88FR1BxJPgHUL5kBXQ+BwQBVZKmJmJiu3MTUIGzxJjDr4XVnK5uhWJxcP+I
1XMml4ST2bOOMvOtEpnnk3VtQMLSl8W+ukWSFX4xhukOHigcrke1F1OX4FUpnmMJ
u62TIqmQOmSpHuG5zYZb3CZicaNYWPs0ADxCR89dWCkm+NRjL22oHFeLnu5I3tD2
bXo8BrbmvHOedz8axdg2OPS5Ghcyj6q/Iu2rmsW/tC6mbUQQGr2Yan04KD+rhQpN
BRIEvV8gNJpNMYJYkKeXAvlfqrsxbGxZ3R/stMR+T1GYMvB51ubV6Pa8ZGUNgJYH
MEMcYbzum/ZmRLdraSzNqEh3HFgbj7+lH9E/uwkKP9omd2obtGPjL3wxkF0Jw5wf
l7PZegRuZN4mqfffp2OLbdT6xlfuC3PlaaR/yBNMpwAN57J9SqpHhj+mvxl82fN+
/qesTZw5eatJ/ZbXRVUVDncpsfvp9FV/SSqqcN7lXxuEafQciSmJFkxEHDj3HEPN
No8zawR9VShY0Tu4OoXZGgr1lFmhW5XwW/a8rt+lp53Sdw3S24CWdPghlmrPeJTp
0wY3PEH8oqar/JQugSKdLaeSQjmcFKjUMyoFU1lBpiu4Li/RAjefD5TN7zuBy+fP
uK6X0Airm+46qBQUdz69peHDLxAREEkWVnnxCAshlXkcSfxnUU2Oq4rKUCix7Chi
kNnCxYNUjVGOleWMJ/L1gxJdivLVj3gNhmCi9LjCvhvNFn6sAC2qyVebponfwEJx
0bt5Cq8EyBzxI48v2I8P7vjpsZt7vEEHUW/u7PVkyjCyYNqFz03HXt2Rcb7VlFkb
HTQIikqzxU1zIiHkR1NRLGOmJlSBrmQMGgzCDr1ksFMVjYNDy8yK1t1BprZVQN/G
aYHaA01DLuWDj3+Ki4FWtUmyvvV2RrTwqJidBVPukx3yJawJqadJOCPV1wonenyV
Xa1zpM6mvmTpVa27o2Ha8ALpjWa6GYpG0zX8yAulhU7DXSX2Xn8z7dGvt4AVPbgo
6FfTAVOwsav+frLa9zoAuMfM0Pg7Zn9PSFvp0lb2heeEUpliVWGorctwk24exAYu
uMOEkbr4vUiIOySGEasrZRqmtFknMszsPyVHQn4BXvjABfllyWMBYzhD5H4Qz9JH
wbLOjg8XFbHtY8mz5LwlKs+VO/AlubWzSsciM2raUWlLNda1LksvZksUXmpALANw
uOg8fPi2XRorMuYwKFYdl0AmN2l4AtIIGMIP2ED2g7KpWPJ+GxYw7jWmzweXtP/K
U5UUDcM4P83VD0dMcqQe1FR6aBwy++M+aTn6Rasv9jN0a43SHOheww5JXDggOe+9
ME+jIyfHX4CYzMzDeJRF6rV5rZJWXTngvp1I3AQ+hYirDqLPLsmhk/u+Tmcwiccl
NFxIngAGO2ptgIwy9xOIqWkCZpqWRRDFAtAhEOKzM9uob336GhIiS0FjMgI+1DDZ
iiDMaxlF78l2DQhGOEphA3bDm0XPJ0MZvxiPe5uhePGeNH5E72E/0BE9CbNY6UMj
q+w2SaF0swXX0d4LwhdrUDPauY4JGHLjDDRtPGsMF6YKkTG3D4fZ7BTszjQB0X1i
MFYDE2kE09AKa9fEw6Baz7oS8A+kVAjjq//BXZv/WpCJPta/ryHetbLI+V+s6Ej/
ijB4+2yGvhFxOjjMw7spYrZVV6epENp4E59+GR+QHpMk7xeJDVPvVapbtWOepTqk
i5F4qcgd4tA8Bf3SlZda0P//jS77zuaajB0U3p5hj2NZhCmWeHJo1wkLOT7Q/bVQ
IY3RClu6O21fRqDMJSQKlONJgtwHZSu8zQsreCquxdjo5Do5zJck1hHdHBXKvQsu
daOmGucFy+VUOZa2bMeFcL8CCQ02gi1y2w8x5fTZFx2UXfbBQz2pT19kyf0yBULR
GeLv6HM+UJVX9GMMsKyHwrkgbD3BaR30iTBAoCfLhzz+qON4MZ2AaUJeiXVANVbl
LS/wg9ZS5MH23IiUXg0heUBIZS11L6YmZmO+UL07b35zim3SspKTTGryToGkuQvQ
FB0hM84WC50OoPha+phfxCAG8PzouWbI+QRXbVLyxL+XbmrTw2UaVuS1WQWzD/Gl
1ZBkPRSOu8tTT8kkKSGoWVwhqNJOkpY7knCincCRWHVu6OzxolxF3LcnjRerkOE6
KAQN0cMWD1DOY8nlasANYthr4GC5Y1UtDw/cPugp0UvUseENs27UgrdL4iG7VcGF
tv6jRQaBdDlzptrqoWmnz+vsMWxL+8ZaJeBlP8dY7kIF4NSKorB8Vg1BtsTw0uo4
k1XsrSTYjqUgrltAfucoZQQBOYf/e/VMQfN5SzFmZXul8d9Gj8A92uyPZxIqfi09
1Qw79k35Vx+isve9+ZhbUrdEv2mJBEnQpvvyJr4kC1++sK9XlQonyWaIg8zbmZ2v
FA2+KdT7mKrgyqoyITqVGPqAG17SmlflXztTSKAhuZWDbnLHCdxIm2hc/WnMew05
76G8VLgu31yaf2LTPyTVdYZHS1CV4MEAcbGu1whySLcjjOXQ3kRpN8U9XuW2qEeJ
SL3cUsmIGGlVgkVQandXpJCapzmDVrl9GW2clA7wfgAWOeVeZMPumVlOHLvXPXhS
/VySpeDzjz/aW2ywdLTKcVX1ukXNyNahycbwPLXSR9afOLPBaDLRTwiQ6MHuFhX4
+5Pzle81VXBva6HJxNZ/7IxbgsYy16IQYfqhjj2eEOVw87AHMmqRrN1jgeKNjo9T
oWmhJnCTC9WtGxsktBDLq1upZb/2aJoyvbYBsnOJzJ3DtzBN02aXE9Ls9XGhzT0R
5sJaHJh9KNIzjCANGkRZF69RcY4MqPXs/umELagJLILdjKnXQAsmwoWylu+hQ8au
u1Ah0pWPlNucA9EM4kGfLIa4SVOdt9sN26Br91mtkD/GUlH40tJD8CSFI/i2mwvP
RW5vJiaZwZxDKyqc55V+NEkqFvTTRvSX9XjWTzIAFJYAxB3STMjKBWdcyy9Cmecn
NYQJrHmX9kcSaDhRYpuOfnlZf27CBpCfH7Z30IYH5I+0eM7rTuZzYG4PwTDj3Fbc
EOl1FSZfF5cIddwj2bLoEmPSEBtCxu1+dQIlrnny7LUOyySrW31ClAPTURbaobgW
N6ZzTXHaP+Wq+TdaRaaY4TcpK7z0YtYpR0NZMmVlRHEtZLGiNkecpcNmjYN/5U+l
N62TGJ93HTvx5Gbq1eqfw9nGdsnq02y5cEaW93Za16YfPjEbF07R6bJwINyZoCdm
sGhC9vudKjo6gIXp8A/9vxU9i2lhd4/dAYFDdIEh+cvZgIQE4wB+FLJLUYUtOf2l
Dd4Ff6rfe4fJ4iPtEk6QRsyKEuXpNf9FQv/+crs3ejQPbqkwvVqPwllvljubC1Im
AcWwrm1x2av3ps5mk8ISzJ6pAwp/XqqhbeTHO/0xZoSV5vuCox+wj46ffpUFkzZu
JhWd1ZIJf+GfWt6EDcmm7zbv+VyNotWufRvWyl6HzRz2BbMXe7zlvF/6g3BJmGTs
mqRFVlRKTMOULcg5I7pftnz6v451l4eKuckljUpq95uhLRF9xBEGzzcWUQXi5jZW
tdaDtoebCLlV/qL9MqhfKtw+cTyJSFSMRXcx9amDVfBmDcc9DHR1zUAJ6FaAtnWu
Z7umAcCj3dz5fiwEhQYgonl97VwTC+wFO2CLWCESV+c6tVZOICBUVh+tKlsmof91
Ea6bjsw0+31seakMfbELbq2/Ldwo/fzxnwWgoiJhx3QMtIIcxaY8jzirGQYEzr0U
ZCv8crmT43cgKhoKoSQoAcwZGsJNTcmEtMxz5QhfKiQqFGiye8PzbRD6ljsBaFLV
lJN3ZDR+00VI0i0MneNJW27U78QyDaXSmkvY9DFRv+YJYzUOxgzllA1zvpCREYV9
PsMgg/JD/5GN+r+6bXINFIkvvvIcVbv4GvCZbj1nfedcc9n5hAMdzP/cGmPCHVJD
stZaKK3sQf41uruFP7mPe9OEmG2CjQgUtw4QCSZzrlYRMjBE/0mskCmYFl9OzpMP
NKPLLoQYxU0Q5CPygkroRfAIfpEVLJNkseMgc45LQHXcw10NAVC64HhNfsK/5T2p
ZhIIhb1x0I6HSYC6/8AXK/YjtdveZMTvz+0FbNkhx47Q36VlRzGJ1IjxkLqc17Kc
HjHp6K2VDeuGGBTxe6ghST4JxF9WWcfHadi0w8IPLiRAuPlLKV6lNnBiv8Gp1C+j
DkOICBz4S65wElwSSWtI50sA/GOAYD6l7FuIhoUtUJsaZ+UVG2JCKmqdJwF26QUx
bP0gpUzqhgCNwxR5WiNa2gEPmpED2d8b/ojdfJZ5PnpnZJpK0PVxzzPzmvJMXj5l
J4ODjGoCryjQsMKHLXUus23/3wEEK2H1FjwOQHl25mfVKxw83ySyYXiMJlsY3yai
FB43CKNgkt4Is8Zh+3rJuvBeoqP63tbZyh5sdGzRyS4L15EZXNe4SXuymoemCgeb
CCyUNqorkux4isJSa8SOrFUDDpiPhhbfbFnc5ws6oKqY4NyenFMn47NDqtxT60jh
Rt4Bk+hQieOecCpHTl+ewkfSF4czNuhUyq0dnS3YGTE44TWxkPXtVkZ0FSw4krZO
Xn2AHXr7hURxRKymov7GnPJDW08wq/90La+swWt+pl/jSMLFZIdvR2eC0x/w997b
WI1hoOKYVq3lA7eIai/TybNbgRprIyGZKzQLTp2+W1TJ5nevIFUB2TSuhhjmYJZd
s8esZ/ChDqgSlB7rJTL0UhBebtUOzb5alLUcgzoZPCPMfCox0mGThsgiij1Ebv9q
eBISozSA4YHymbtK55StCv5OG2rogQAVZsl042aKLLGfHsUC7mLzMU9wRQrOktAD
ilkpl5T5+WQ492VZiFuk1OnKT3SpjXOYke332ymtVJprIsAktbxSG8ynlKxG8hqX
9pYNYvVk6xFokZu2ioQs7XlaZEO5m+Gji08Qv/AeYUUjzuIXff66sFjG4k2Ulomk
JlrLb2q3PeHxuxKybJgeEag7V0dmP56bWA30pABK9y+tLgZbxYGzkoo9W6O0D4wK
Kq4SGXFOl5YkUXMigUEcEUtofMEx0H5phb7oky6GLyOkaqSkxkeJ8WErMLRiuiWW
MRgZq6yieX7ZsDFX+TAhsQsxNvZZFphxqbtsbinUjtb5U0ObZKspeVZNQ3LAXcn4
xN1z2lX4TDpQJ3YeLPfhqznj8x+mWDK1AXGp7HYnpesYAACA3wD6izv3Q4jvyzVc
iv8psYqfW6xUtdt6ZTfRxsvD2uR3ns7B6V3k0/+WH91es6p+eko/NvZBclgHXu9Y
vTleXvkPDx0tKy0C189RjnS7dmN5wny2IoUyoGaFEZihggONrQKUuan9wyWhf5xp
OCe5pUa2VT1a6wUBl0CfF47aKWkuLj8EN0LeAsalBw7wIPXzC+1JS27QV8C04WPf
h9LcXbexxlxB0KHj62hNrna5IzVwn9HKk12h3sLo2vWDcketOjtHc39UbB4eu9q1
wyy02kqhKnWMr/+JiR8Chv0pKc8ZEoolhuY7gqhdGRbr3sAfOrkkwN1r4yCqSQGT
pa9GKT+ux4nqNtYxjLsOmWl6Qbpp0pwyEy2UKwS/4SssLL2QQzBYvThCuftro+2r
Lxe0x78aNZ/Su6/9bN0iXgnk5R7mrdZNNyQ8LpG2sIlcMYdpIWXTRt5hxCi8YVrU
aqNpVHDXY8tBxHagLCXphip31HxXNT0IetB7ufFVhH1LS1kR2nN4YgcZN6/k5fcY
ERAgj/pzfhIEozDsVzPLlsT0x/z1Z6pr/e6App69zPn7vg03mnSJuxlgC5yd/Xn1
YTbKYUFEhehyXyXNStjogSuRgYfjxsmtEYtuzfdaekI19/CeqjKGz/Do79mlVzUP
aeBroi9Gf25UdcKTK0LtAOicz6mn3PryzAaHRzEk+lVtO1GWyRdDxJwm+J8EUou/
+aokkvaGFZsOcj1LKoAF3ZU+PYFsXR10tucY9AqP3vmUr6pYErTPH0ZY3TnDbkYq
1bjf2g+3C5mD9/CYimnK3F8+ITBNcBP6Iz9r5eq3CvCyrOylbq8EU4/tCCKmO8el
qRVxObE0EQVUxsnJk7ZcDG5curz/QowIKALrogqCcWt98zYzFCmnEI3CPkryMfdN
Dqv0loLuWUDj6Bc7VI+Fqk0Km9mvTUaBBJaIFUJAcad7RLmwpHzR5TM63sTtlMoO
+W66aBtlGC1nDYQ5iICWLxl1DgIaE+d/1wQ/R0J1hoC8+H7Klm22hm6JCj1WLJcW
X82L2dfH+8wzHwxf/bUeQqoJ7rtS15ZRu/+uJugCvpCFqdI3cbDHhuIUxnsvb2+R
syZTpKILu3+ypMnAcAujMatQaCKwFOlmktszdFpo+wIuPMgclJGVzBww7MB4i3lp
K9ESq+SKb8Xt7MjbXSqNeDdh7V9dFM5KE9Cl2eUueCR3XgQHMLfJ2/mZl+mXi2rH
yEIxTX/9qNiDovMxAlDwGlMVh00r4Lk/A8H86y1CFIbycwJHKfw17lCRHA1eEyg9
N5bNTA/GAoUvyd+4RLw5o22F1F0QIstSRQuhggU9SJj4AWNFGrBpOMdnxsBPz3yQ
VlUMDwAB3fVLpLWhp0AeqTEAcK3oBDUOjtbJmv/CHDUuKdcwVuB1lDHxtYzFmSVi
Ufk3QbuqJsTfEfGrPkSOCyrznKEaGAdBDlJji7kb6PB3daKNhqaSJ+VGLzjc328F
7U0JBQahKnDrfDuI+bsNg0Wec1rXpbo0LjdVmGZaa2wbxqUpzgtnqpB/6LE2Lcjv
Nl/PQD4VIK5vrxn6OXJaNJYSBrRVRbD2A9E033+FsZmVcK7Uv8cdTwXDeqs1yBbd
TFMioqzoW3SBYXHErbAgi0Cr0F099toc8hzR4ZKdyJmCUJleZOgQZPY1o0n7/I7k
OtmbHvbslmV/T1RfdMZZ3Bn/HMY559UNVI4yPO3nGSPpMsAGooXiyHT7mQWgfKNL
hB1lg9ETVs7xSJ0TTQUXIES7KrILOTtsmm09PrdlFQ5i/Foyn8v/Hikk3HT7LvAf
Km12VThM46xssNW7xsux3Dxhc0en8TGmGJFiSGCO5OgwL/PSwihaIpj60amrY49q
N2ckYDORF+5BBKP7ewRhOP9mydxJs5OPVDYrLBfRxeXzxkZm2ErhxKfPx6qfeu/d
MeG/BU/7R2qKW6esJJTLQWbPBUnzaHHC1ZxjuOZqiqqxg6RJXbQ/xE20FeepiQ2u
E8yjA7e4khlCGaRPE0GxQgEF32kj5+RDSMw47Pzb6J40M2d0ayKuRCaVPoQ/JG3Q
GD2WkJDlRQDCVnNTceUh1NUg1Ku9GcVoJQUnzl5BurJXNK9gNKalKaM5bopNNIn9
3yWdTPd282ckEB6dezpUUtAaHEOsIK2N8ocZz77lA9Glynnlaf9zCvKL/Iu0EeX4
c3epz8SlGhoQfVaTWVQf3bVKYhZxIX4twI/fpbPmqiHi/y6KPT0x99CWSXVR0WzV
IyBqjH9biG0z0Ju++R8NzicCy8G7wLZetaNN1CsdRtO7zKZ/KguiGPdsvQhDfKl2
qkWo7sylKoILNhC69Y7Z3DaKlTFePZvidwRJt05fMkBZhaE7ZOR9RSMejAYyEacC
QHssnqlwmHAytzq8WuxxtG/cXTzdR8xCN/H53/qzf6TJh3c/IpcqbHDRWQ2k/osh
ynzBI6wCRxZ0LNLt0PKhPejSodvDtDwmflTdM9YCZrYQMr0Y6Gu50UZ9ubWk0FHR
/2EJgn2NRqoUCpwrjl81xJowuLPEhD6SzNWZHb9nIKzrkbDdch5UL6c84gUUTqoz
OPhDNBjKV1I2gPTGPsb2IeasagQf/6gtlI/umr2MZrFgLOHWdFWHdIBtD/xBcqGY
fLEt3NCptg/c5N6Tz5KzD0FUOvHpgVMjCp6TVWP7FxhvoXAFeQqjN0AWvNxQbkV3
h3Dy2g+4qFANZWNpoZ4pohZNDYBqtOVimTzU+RkT8Z/e8S/hkQwRv2iXziSoRjR8
itDCUaALsRqoiVFyLVwHp/1P73rSE4wyP1uej2+pVNRT/az3m/IK4dgsezKp85PA
AHjcFHyrVs01FUwhRspH2HoBSjSVrWGgzUOALiTDAB5H7Nq8oG3nE4+1aE9UPcR1
d1si/4qYiAZ+SGVGezS+l6P/X3ZhpIgy5u0kvw+NPzM47jqmDTHJLuVZ+Xyec7jA
tv5nQ6/kSBA6iGF2ztMlmUClXxpOzsuTF7YFFaGJLrs41dKFa0Moqp1YwmSWtD6X
ygKRBi72Y9n7ScdYfRH49OHaJP8Y+ULczg65cWkxAWwc2LUnVh3FEcn9AmNoE+1n
mFThfz6UdOT5SEbqjFDQH7VxFiqlMZDPbLgm0gkkUytEeiiWO4kSrpNt9yMGFfTB
itWtr8cFB7yQE6Di1mlP1OjpiO/pzchT4PX6xEJsae+Giu7JPxlCR5gghMwahaSw
QzL7V37D6Ax/C0Yy8dt9FkDD/7ijj4ZdGQ7GTyB0GizpHRnfZEUDpJow6tOfW474
XMniF6UhNOn1OsMM08WxE54IJVKzFvKjiu9aVRgv1HX+LneDQx2I4aJYhBYDbVEo
B/0k6AEWqr1995Uf/BZnYomhsPXiw8NfUFGDbhb/9utmil3fP+xzNR5Oa+JRaz/M
k5p5sUjT4ToXzDUvf/rupjt01xQwcfiNOLrHw6xivQDCCiqGYTI8f5Wr0tjumsh0
J0cafsEcSfWNQS4DekBFQf+A3heLxROTg1Xqqbv3MzDFxfEd35PlyUFxcHkVrJ27
DxSnF33ybXqxSgz/VPlu8tYn6NaY86KZbFhknDO6+IbsELLwDS5RzZG70Qi2xFBH
QmTiyYQdyGJH1J4peQG2ogpTZ0pleaQUxqcvbFk64epLDdMYlA7t5wT8H/JWgsUN
idku2tFFNJ8DYUViY3798D6hsnePsY63sSAgUhRAkYTcfO0BM2Z+Ogaw+aGsjJAj
c+WgVVPVnoOTCOUngq92pN0lK8lA8Aj19NQWANSQCRNtJi74Z2fCZFLUslGINTBe
nsI57H1cX6b+YsXI0Lq/OprDVIK87komCsQupqbQe37MyMd0BoA5MhoQmvpn2mK9
CTIeyVdJ0YWq+/iKrV13xaf7brj/ynekvAwhI/CHSRw1kS+tXNaV/Da+C+q4egcL
sX9+zcsty6HsQdHvYz/tteatDfrqO+WUiw+v9Rl8rT8O3vJb/D0VIH6Y3nfLBYzL
Q8j0SYfqqtqqyRIdEqEQIzayNvl6ppVUkr/M5bjuhlZupemUmEAnnKumt5w3zEEe
m81dfChiiEDyPljzTk/Y2Azc25gnz0VvnmtPdkzix01YUiy3eIRVL2aZm88I+aeQ
t8nV3MPR77/Fhl7uz0VCBbRSzvYKOjmrsG9QmLaQjSZsk3sIJfbuHNxEKT0tVIQI
kKRy+9uSybw9PM0FiNWBUi5mzCQ8sm4x6UUTol2QakiCN0xk2eWcVLFRcYupeWnV
H5YofjifezNEC948Bhn1ISdyGoadSYUTdHDewnzAZHAqofuTz7Mk6FrDYZ/Wb3qQ
oQ78L9ICmUtmqVqM3piYhlNsPd+N69x05eSiuhWuz/vkxGnCCA6JEIAHle6K9k5L
Rkbt+MlqFKEeqwTjWmhIyQFyPvjiXQHie7OmDziH6+AyOMZgHambDgdxzEbS98af
KqHdNL0K9Btm0N7f3b49fhfT2TSXdPyW2vsMXEV2m41BqEW98Yg/J31Hofogl/Zc
6IViI3Qy+6/Bh8hLTcRWDg3w2LkWHIhRvyeOltZTuQIV+7Z1pPTKULynuGNMMl3a
KXcUObKwmNSq7cPAypSZHKHIUQUXmjOxChkt16nYmHFarzv4ANH6nmyexpOSFYH6
bGzisLB09C4hgJPUmhdB2o7hkZ9PDm7u6ZM6bBnDq4QPjruJI4rg07kq6sGsvnjm
8yjsVo3KueUMAkHX/vL5Iqktu/ZGzlk0iITR04VlBgHKoDkhLYOJjws0W87dysLc
+SQaaBxgddY2qTxrkuOzQ+SfIaCbqjhOIeyNFzi03u2xgf7uJrZ0TB8mbM/PDYyB
XDVU2JKGiO7wKipCMMaHvma/z9DR2mirpSXRmGZfYIv7M++duw6ftNsKyyVPJKwQ
SX1EbUTphxWEFhq4bm1xM/nmpfOCS9h8ycDWKy8IS3Zu7eUwkhtdpSXqkTPXCkVU
v7tsGT/QgURgC/oNPwM1m0rFiVSQ9dEq8w77yqx8O1+LERrLdngZT+SY3FT8r3XT
dYZ8Qm0uLTy9aV9T5+b/r4Ji79HsN4MexRfNrD3MhN5j1TsZDatp0vhJBn0rEaEm
vTaYFOOzwTRM4aKwD8Mhos5S79QqJ6SbEuJki3DYwV3aRnJuloergQUatB9z+VBD
2/d9IMFd6MWFclzATwfS82/oQu4dNCbdKmvh5pO1SD2lFDxWJ2rzbKTfQ2SSR3E3
FFThrtUE6eq5qt4+jwnYUyaQ/OgT2E5bWKeyYXD3O3qOHlQ0CDgUvs73ZjgZtuTy
TU7zAJcfcGcky26HnDWt2NBQUcfsRAUErIJM9gsPCNGDG6G2INhCsiK60Ky9Aj2y
zvx8lxDGRXIGFfubrzZTbrLX1cVXC787ESfyqRRkDMI50C8ALa8FaZb+ZmCN9jiZ
KJsaOSXNvyjR0G4RBge9H+uneOhNJkfLCmpgvWwu9MEAjiRDQnkWNaOo3H0RKfqb
ngOOvrthjQvire2EPYOBISi298IuaozmaFrb0UBPeBsuDviRWBvm0PFhLjyRPgUV
edbdNiqpKy/9wjcgPDDUr0/w5grpdTkBINC6SLG13akITY1QZiA5743HMi+Sgvdo
IaQB2F2OG+vQaJIBJylAyHWtgrU/uPvFeHC8VG0zdrqlqOlD/MHMDzhqfxbRdjD4
aUN/ZDHFEWbyBnZQYyIx6u0adWietr0QTIbC+tT+TtAF6jPNGKrfJC2xt12UsH8m
8PS2XjCbMl2WvvZu9OJWo8iIFp36vEICrPvhydgjW10EAjb4D8ameNfuVT3qN4k8
XkZ3iRPfRdqC68EkR8+EbprKai7nv4XcqhTlv4HyifCXk+FhYR80xk14Ln5APOSS
eMOo2zlXb2Gms1R0B8ruGlZYa2gCwp0JF3VIHG054a8zOja84AkHPQkPW0+JweJD
SHEgDCCYrbdkauTyVtqpdPMHk9fHLM0XXkSlDk+nmHEiVWKruljXenM02+CPvNou
nWTQy+5+yxi1tLpa4VHVBAbPL7D+tcPv191Ad/uTfrT5RQhXzrGEp0TvIQe1j/tx
b7E55rqlO1hkAER1c2x7v3B04CMLIeeOsHEk+WfhV7f7J8tMr9yPKTC6Y31YmZeo
aszZ/PHMTnVIvdwebcVwAPsHD4FVi63JkyU2cnDwChVpRIQLGKvtHrs4u009Didh
uFel39FRns/epmmINadVR4ZZct96TndCuODhzLpYjxqPJ46Ne5sKrShl7zUW5sZM
Hxq+hmuwHeu7ux/uRN6P5Mhm8My2IzJyodzNpmBXt95rBDmv1+f9IMjQIx846iEk
8BtUDHH/uZMhE02SbCmxRw1FErcV457ufDmndjwmws+So/pe95cZ2hKQcJgfG4NW
l9WW1At5l7UxqeRlI3ZJECuryk5en2yIB0SRRZkEbMzid9iMrMg2Ngvk6U/y6Bzy
nR0KivQfqSvnrfydwFRdtwghkvRfanedADFd/gJqTC5z0UivYBIixUmbqbXbmqm7
W1Wl1nsMUTyroRVA+qmRX6rr0k/ReXnGEDU9NbRqPny5AcoSOwfPT5sQhAmZdrdF
KIk6Cfk/1CfU8jXRkajYXtRJwM7ZDETlEpzWhsIVjzx91P7SctaPSe4uBBIQlDCX
q5LQbhpbkHr1LImi+Cg54IhqL2BSOYXYPnlSbJEf/4wxscKRoaM1xk4WtJA5cW4G
keQh/R6lcXmlsxjLDAEt98LSPvf3/7YbEQ9ZBKQLcYM8V1D+WA4iUOBws99vuwbr
NXjUNAkef9NZuGcf7rvy1wLLjoLRnHTIp//qal7ltD6b+kQ2QHe7+qLdki9BD4le
aTAHoRustCfx2aa2zJzqZusPUFai0aD4UYmVaxY8f2XYch7Kz9Qy2qalZ4YKptBL
9Fh4IL7cqB0Z2pgLcmSLdHVRhl9xYab8egkyyy448XEqS36i6U0FeHm/EwhA2Qvs
IRfy+/e1aQHWvwNOvNwScmAgN53v7ovkJU9hWSDwcwLZh/q/8XmWHAoDFSalE/jc
m3EAs6maEWZkYxfFATw3ABo3TOnD9I13eO6JaPTGFhN9zt7SKIHd+7BWJgavCydD
ZhWE2MUv31bov6IWc1PV6Xc2iHOgh9dJHVRnV4SFz30uf8yWm/2wqvWzxSlyA2Xb
O9F8liebIDu1dsAQaWq5lckE0R2mQjYTnLTeciNhai4ZF6oadPnOPoO2gIh0Mk9d
HcitqcNyYBenmJn3U367YzU2EPObCN4RJCUwuCQWQPIdHH8WxEM5onJS4/jaep4t
ZikP+agzGzyuRmfDeJkpcEj2v4nVU9Uzds7ThdqVdJXyptTGQ+JgZxxvsdnH+F/u
XusyDoSXykAYp8KzUKQc1xHz8Zsthcrx0lCJpqzj7vFc3oxWjV/nKlNEmDVcitnT
Xt3q3J2PLCQU/pHDXvmuh7dvy/M8g4Sc3+ZdUJVCYtm4EynWw4cjkbc/LqQf9MFt
ycFPdKyYqslVKIaTr7qedeuFOqTp2HE1FTOxKS/WzwGYTIfkuYd4dyf9bnpWf87z
D6X62mkppIXlRfZzwTyW1qJXcpaDUNtP3yalSj7LtbGQUQR1iEpkhEBmzqd3Hove
qUp9+VzkmkJ/6jCMCQuRDqrICu1TbyjiSkZo4XsFsfc4CAmInvkgyJE2jCqRAyOI
3tckZ9Qw6jneEzESHQsxAdHbxk1rkakEIMMnjKdVW8G5xbJv7b/Y4TW9uc9JLXhs
oLANin7p6NXvIrYLWBx4YsWVJvTpL+5WirYTJ4+KQMSbJCWZSnY9i6h1tMne+Rya
K8FNuen/U2xaVvF6o8k5lLeStAqhJ59qwJC7PXM7OxXIu7Al+V4zQE/6JM3qcz7f
W4PM+btEgE1hcqgODvoMl+L4zxE9W88KtKVLFJzo2dAFR2/Fc6b8yMtZmKi9cbx5
r8WmCGaJVom+TIZ58q1x4nPcYDj24TPpq1zl4Xa5XR6sUFJhpl8RWzZPApPb7gI1
mrRNnO4cJUq+yS3exuieQ29tgRPFQ/3VastXBxW7mdq4LDKEsQnTNxeXS6IDTJgq
m+rOlKUs6woXeTEZCJ2QshA1CWANYwiFUhhs//a87KuD2IlkuJ7hvRnUINYpHpq0
aHkryAird10e/MLhROPuSFVUWM9SXF8FOS+TW3KLD9u0QOeBqyGsNy06XzcDZiiD
BAdy9+BxsIUii/XMSFY3VLkCMoQYrOW5EyaqEXlo5LDf6K6NpVYTp2e1KZOAEvPA
2ZC4/epjLoku/BgyzYuyCOxaqBERGoIMLBWUaHaXTa6UHqKR3fRncNCbv7K3b1/W
zPlt7cTQ8Ytdn7zIRCrVILEzNbohYdtZE+muX9uIDYhTmTyd+pxaJXAGldD/vH63
C2Yh4Xe1XYG4Y0nyDJnMJ18Ji62GfWQoKszCRiWYn28/ENZFKDUgoX4CWhtw1O/c
aTY9pVPZkBQX6HegTbovZ3uOUd/rBAoXzx7kuwk6uuHrprZyEemY6GCLOpfRhjwM
NbgU76mSPYis0TZkOZQ1pwKtQn74gjAbTx/4EE0/bHRzbz40iN5DLNYJAvyF4eOr
xM4FE6vhdjS6D/7ClKXAy+6cRiYICGPUPiHWkjrmWUJa2Hu6xyzz+NcVL1LJSXi5
LqXp8scQqBsEuaIyP0fxMxxuCZMq+ix87Vs4cnm87/aRPlZM1m6Oclr0d1T1Wenb
gUraRWGMDEPOhqZQPzRw/cQ3/rC6C1XblzhpGxXP2ENRNoCCQ0x8cbsz7SXZ2Orj
PCXGvqnwMUhBe+/63DQqMcXGBCENJtbixhYA64ZrH6eqbuLvFgCrniN/aLmVz/hX
vju+FgmrwA7ZEbSFmbiTZ6zSn++kHeGhmJOasGlJTzmU2ADIvGRT0Fwsjxl3EhgO
PigacElYjfDnvAzxtx+gqwNjdqy7SHseyrnd0Fch0cvxFBGKPToKFB+1eMZ8KCXj
4gFppUA/3f/BxLzeOdTHybZ6SCWQUKaTV0pV9MTCc52nQJXmbPnW8QtlghRYs8ml
viDvKgfBqc391HjoD16iuT20QOeRiTvFcWUtSKYnT4OGx2gxJ9do+tkuatSZXXrp
yRL+FxHYsais0I0fIUHQn/YH1GBs4fj91ybrxVqCcO88n49yD7kAlvZEFcl8qShf
CpaSS0nuHdKBo0aV0W8Z/gToKKI+I5xW4eqYoqXmTvY23zb6C9Vb22DwrMxPJXra
vUXKhL6X203FZGLycMY1bV522cwvWiZHLeS9qeQ0/DvVvxCDXb3R2PcC5qU89QFS
WN6q8FO4vQg3tAmXn3hvlB7v1j+age5q1pRKL0agmZK+w3f6Td8SvZS0KwWFOmaS
vCDp2QUc7JBwDE5TgPb1JDfu/BHeXJ5+QVOs95+kWXZvS+Wur6GUieUDXV8btV1K
sl/bILtMhoGkBK7MNcnxsnHwZvK5A/x4UuPO4muyWd2O81CUa+zENclCXxUcL331
TEMBgb2AktKhnGWfrf5Bd0Lbl9Ff6IjpjMhB59RcfBwJbOCeUv2lxjxjsm28C1ZS
CTrUa0enxPM9OIaTS8cZyjKsoSSgg6/bv78Zo+xKNeVbz3j2GCnFW5cxXdruFKlm
MaV6E9Z9dlbdi17Y1yLtX9peL7JYrAaOQg0bxYJnq0ris4LaYvQQByluOUq97yKh
Ir/gWDQGGS+TPzIWImMVy82ZazxyRCOEc7Cv5zmzCBB5uZTKRyBzQ8xXrxhrjX7C
WvKXWjLGDCr5sIR36k3iOK9E066VlSYOXfZ5gvumsRPHmf8WRFAN3P3u8K2VJ584
PL3AeLP+Qes7VSwUX2YG31Vlzt9W0WOtNRFD9KvS9ZLAu6TT6yP6Lyum4FpoCf41
Lmo3DPJnVOr5gWz5uMA7PwYhE8BtYvW5mXlP+t1FhL2Yffbjt6GNvdHWQTplQJOA
62lZUUUhnMkBYFss9Xescq7Lo+SEmV3zjv4urxHoWJXMOCFN0aaWPxACOoVybcPY
NcXgIjgr3+jCSvHAivcmKtxXXpVnojJzlBFvsNqqT4Lp4ywfEsREjmxSGXEZ5AOJ
Wc8TmblMtvN2/dp6R6y61hzoQaV0SmwZKwKYZh+Rvd6SWlfXCZ6EvXr6Q/YhsfGe
LnC8LEVVEjICbnDnjA42VaLhpmuTgjTbXDmGlXBgh6S/LPQzx1HVe88zQ6AQ2Ag5
ULr41Sh4yXTNUZwtMwrOkbCHlZET9x5UHVZqmlDU5ZBowhVeYBVGhjAtN+oR09a4
qQloX5mRh8uttNbMt14B2eyh/45owOpjlDDlM1ew20vOcb6O7hXmJTTtf0PYQxdf
ElXjtyf4RwHTpEfY7hrLj4ZXsLfgTXmoUm63wsn3BCrCw0yyISliD5xKcIKOdt4E
lFkCt2yMOGlUIAJCWuRfYxJEvf8A5ZYPk78p788joRtRhEHlsRymAS+F/kL3Yqdu
RKggT5/HHF2qRKPYgQKAGcI+Q7VjAs4YxZlTgwuJYFFrt6mBgV1hBpkQiyE4qwM6
PUpmwPaZQtGHslLw5UctA8ybFq4QbaoMur7Zkhij1ojqozVlTxIczgHTmnIbubwe
VSsk61boeKD+9us9uS5xSv3qKF+7l1hinTZf06UoQ5urJL77hb8pWfq47t9+8rZs
pPz8YbRtaZd2MDb4oKjRNCaRN417XlYZPMx/Xv06oxKx2MyLGBrqYnDy1JYeL2wy
fZ+cHVDwUP2YI7OmuNwvcAYCsKNKd4kBF/zVofT6BmIcRO0KZgRUbtoOEM4LPG92
VHXK0xH+BooR03ueDltOxZgstFGhxMYEPb2rzUWkrrstub+bD9eD1ihFzvcslS7m
sZMIYlrxEhEncJmA7eXtZrESBYVymAPdgKXQehQFxewi1CN46f0cEso7Hlea/WG9
f3anP54qth9XZ5KPpOTHrlBwmtzi7tzz9A2hbyXhyJZo+xUc4DPpUStqBSlgyRbc
uYqS7BVfgSXXFoD/dqJUAQHDR+ycL4RXqgcCUNyoWjJ+vDyUS5Q6rtFBydQV5T2o
P9SZbaKLKhIxy72OJ8nHWDBg1dSyaHN2ygvpHcuRHw2P4zEwdreS8lKCIcnckMbw
Bzl4Wv6RZhWc6E6UP8ImZuHCEfBlaUp9ccQTHI6VOLuse/oswD/EiW9d/O7csrkG
lnhewugVDZt+mZ4zpQm1qcxO8RrQDHEru1A4lEdRdjM0o8H/wip7Lv6xszYABuG1
BxKlFlCR+Hh3a+UIseDuXV+ukIriiq3WIrJ0UhEGJAYK87Blq6yfLj3w3m0MGvoE
Bjcu/+Ae4AdiL97xvBn18n9PgAbhw9/NdkmtzDKQWL38n6Cx8rEoGXhNY1X+kAXK
OZKxRzQYT4LE/s8fluBxFy0vDnCy0jjIIrkKCW0JfA7Btpj5AWE/WcNzEk9gLx3H
krf29x7nrTFmaDzw6V8J6HCjENV2DjmlBBNJ8DEn0ZhKo1K4heOE2rYpy4mm3b8S
vOEUXIbO0rwuXpoHGQm5EcpvTyJPCsmnyRDPZj2k+64ehkEMfAXZR+mqWujIuMJI
nMSQL4Nuoic9nz7lawqqqXi/ZRUkXD2jP8JZMLNmLGxTKcTkeOO/AKBv8T1vNlYh
wDQuw0t31q9tKiPymmrbRpPRlKQYlFjaRaxh4fHET5IaR5CJvEAcxxeG17bdloo5
jsqqLWCD8o3jzrmhlzxfgEwj67rJQzNmNUF4ExzEOt3SZH/gCTRZJLyuLl3Bt1JA
+YCj609KCrYf4kFOU1G1romVO0xawPeCUuFbCGAsJIo8j1IqAfKJ2JaAiQXAaJum
mSIa9aITi1zLHK3QNNmjwdwR0C3rpTQRkiEwl9dHfUPwHJzBxlF5oN7YGCVx4mJj
4d6GGkUldY6MpcjVzEU4zAv4OKlgf3k6QJomDSJW/murmjwIwzxJOTQm8pKsvecJ
BkTyLPgfPWKWq4mqDP7ixGsKqT5nqQ08HeDwzKhunszhpF4b5ffhUuQBSqTUgDg1
U0UgZEiudf8+3Sq9/pM4cMuKPz+hIByujFQUe8UX0RZEniujs/fVQtBJZHHhwZo3
00KFWInZgxS1pVY84UHIaYzg2+2dd2MVKJ2DS7uZe95InH+ZwXiMXq0yWKQ8QIp/
A71KtIQ5NwDPfsr2u94Mr9ZF8ZZI1Fi/2TEC9RzSlLGiKjNp5b/Ie9FJ1GKBcmgJ
IxgoYpw2X2GoGzeiB65gwzlZ3nCKar3aGXtwXsPWDEBNKEV2acdLyWJsEo1Y4Ir2
5hL0c91eAjtnqHPwOsIha33IOJ1zMpEv4PAFftgYUp8xqv4wTw8k3c3taywCiLgo
DJ0LljzPnIlk/iFaSdLrR2reShnqptAElEesRuPNuEMdHqBJ3r364nduAFTTDgWR
Ix+EJrKhiOBB5KZP0ySoPIaeiWMnXBt8DA9pmWp1vhnYTxeOoL9dJmE/TcjQjWYq
J3ALcpxyIhtNVhW3zzWBUNPO+SfcXeHyqBzNYbOoloOEXACoNycg3Mjtufrj0MSq
LSr5an2U4OXtQ0RNKECyfS1Z3F5XvgsvAntxNhBStN0YTM2/gZps8sS8ZrBmWX4p
WjE2ZQChpwO2EwOV8yJkDqrknjg+7fuOtyDbiUxtXUrg5FQrJH1CUISu8/j499kI
gEFzykl1xmggvD0obl1d8XolJ3LVDyZ13axn/7q3JutIaOrXuo9uQdUbpB6uIfT0
mZmUPB9Mw4bx3d7zJ+g2DBqQNOD5H1FEkuw69ZZSeiF35oURZ1Z7Eqm4inOO3qTA
rAEEwf6dAkwnn9vK+L+z2jLTy+UpcizNNwqHILrvd61nLLIpAWzTnI7vqSTPR16I
s/DsYruCa+WpMyJO/Dw78SMC5JnzIFfeOYYBB4NuS/NPUJrEJGKuLNbHwyDirVQW
DmUx+7wnksm2D8ODPgqwnApTcVK6FoqVi0HxQXc4++49TAD6hXyegD6ag2bORK/J
qvfE+GT06JADPQlIaggSDpDCbMYWRpJmD2NEu5eCg2OTAMY4G5klNSyxJce1853D
1q8AM9/RLG1w5wTmOHANzpbVSzVrH5id9wLXYRkjW519aDR9pUDmuycxQwoEiv4R
X54cA4rti/YQjKCwMOmGGzK1kl/VjGz5ouR5if7iV9lqISmgK60g0L9lNxcrzle1
o0e5tTyVgvk53r2ckZ1dRQwS8uBAzx//fgubWy10gHHiFDkJmV4uDw8mx2QQdNjv
ASA4z6UPGv8BW7F6b7Ge18bj5YbQC/b0NXt2wHNxr3GLN7PIuPQQvPIbYnBfuQYR
YJce0rEOHmyWC7tFx2ft+/v68dC2rBARZDR7B5St5dFrCFujwujACT8MHI08o48j
jYFNEa2WnHcw76q5m3WKPFT+jJXf36advCQnGi+1QHgVuOMxL4f2zA+UIuuZHevm
RKBcWfXhgwXe9dRjSCk1LLOk6KnZJTvELSZK6w2Gx9rQ+KomkapvJXCq07wnjwbN
Pk0o6V14AGtQ4NNPpfLM0VTzrm/MwwgEPnml5ss1cv0GDP902XcyHOD3MDOnBYAa
ZIXfP/19LmccJGwNhkxzLpvhPQOIZLXoE2IGJioLQWoRGxhBdQTRAXjmYpgb7gOQ
4lM2ox55WxShJe7Cm4WZyibh0yAR7dwRti7L5Xh8yxmwTbWFvWpXqWvK5/9K1+BK
owl2TKYnO+XjJhJwo51ljvR5Sxpxep4y0m8r+tuHZllXMYfBdAXjTlcFpyfPqr4G
Qgxdd08FCAJuxL4gRi87IZMAYPV1c2Cz+xxSAToHW1YNOGjFQdmqRZltnJB+erKe
w2v+QtKxyjBXVAJ99WfF2YM89NIA48WvDyjF+H7iCNZPop16rJ4qvG9yqDowfa5d
ws0MRHqgkSsrfvIiH9koyYqoJyvpYO2cxNjp5GIKC2tY4FHjmaRGRiiknpChHEfR
GKADLr/t9Bsyj8qPMTDXl0qEG9X6KcKusaZxHUZ9WxxZusTgt16zu/On3KhU0MY1
OjjTZ6ZNIsqw2cNVRzmAYRsj7CYmaG4OiNbk7kYTWOM1bORaEVaxq1dbqRykyV4y
/xtl9GRCGorCv9+x11xBLJQzn+biZ+C0XNNiJGTz4M4PmwJN0L/BHly7lFCy6q2V
Sr29Tg8SREtWT8Haqs52VAU7BbdtzWSRM5gXmyzdyPV8RPsRil0HsAT1Y2xWEBDS
bX/rUI31j8pSjb7dVi8R8cI6JudkWDisO9KFDVDH89BMKUDCEHj9pemtAGK9+SzW
rQdh82pkSLh31gORql/DxS6DyeipPe5LMfebw0aTD+QQgvb5tjQbWxPCBkq1boxQ
Vk0um0sT6rbSvQSC07CmKNrnXNLqYMyX59LDopXEn2uzs0M7XBzCHw7PUNEAR5cm
g21LS1naxYrw46ToVXJA1f8ZJZznRcm9dSvZ84dLT2GpRn5Bi9GHfeFBlEMgVgAO
b8peNqrUw0HGeJYDZ90NcBX8O+sBO4RJaoFkaV0B4QU2XDnwh17x5Se/dAcc9+5w
D+B+zic+f6B9d24DXbpSMysufa4CawXiE6VK6IGt6hsbdAvWQdKrjFgoKt7iEqT5
j4JFEAfDjkKKX77no1J7Sq7q863/UygDV68YCwBf4nWs3PxqTHZ3XSg3SUeC9pyP
g5G6YzM365kNxVZke6CDKh3IpQ7SZuHts+X0fBtof4iMddn3b6yrWra3oegdGk7D
N0Oarm4UJjDJRnbcplAi67+UPjgtSczU+2RgbI8GQpglC66gRRbaWLyU/N3OTNxP
rWesAJCnOhPlhF/l/2GwN5kWumi0usWX4oYnsDcohG7FejXzupo/yRhsFFepvsBm
K9LNqir45B6KXpxiTz0tyDgyv69PcWrno7itS6Ah69/kdalOkl9R/i7bdA3daApz
lG8ZicO3Zs4yiaW+H8rTwNvWihO8GLfN12B7fdvIFNgQFYHUh+fcZj3sVl7C82BK
4GmG4GaqIDH0PtSoeaEAv/EaIYpECRL/Wtk9dwJpymlitoBnbLpCX7gHViyKKwBJ
Fsx5XgOeSaLMBmSnP5yswLxqye1u+8N/vjZi6pkpQGb83aqSGKp8BsE9nSR9K1tJ
I1RsxfK3V0JvPTHub+lzDZA7X3sh4jBsatSrD+YPpKeLLQUp5TmVj9f3wtiZs6fO
qrYznQUgQB2kyhBjdPGA9JdFvl4eubBMlwKNozUxIAf7y6d/ig4i30EbHXoksWNu
25UAvKNcC0mb5yyYBSRCWR8JvLn1YBGiDuLEVlJnNhu/Vj50MzqRXaWW3CXUAmbC
QYHisM+dTY7ZCK+mpuAXd3SputS10bZaMHHWXWBZ7n8GToQzIopjY3W8qfNFYNIh
Y2/O/5AFzfY4RM6PRrSpnE8V56K4MCTHjLIzXc9MAysVzsSvBBosDRN1RzJ5r3er
eaDs9mhJ9hgudDT19gVWDFGiHaL6YQacTJ7YGklAiVTDUtMsDcWWuxm5WWZgQY7Z
QJW5P9dpLnbYr/WieqdjbF0nGtE1MsAlWLZ4o1CJIt+l/Ynmi4OfKcSJWIICVjJV
TwgL9aMck4MBXBU1jX0cUtp4yRgVijKDUBHEnP2+8azBkbQWSsIaeMtJryUyC6l5
ZoowrPhHGSGSBtPngvYGoTGRz51hbsmL42dVw9Gbh32z04K0/LZ1BFYlXxEMuKPR
8UiyKPwJsbnQLa8w/yB5TUWBUR77hADGvqlP4wnVckNDFAOEhmOkDzhD8i3B7LAh
YlCu7dZCEW84KeCcdl0x1jWKVF0gciVIiEGNtkWRfprFzVwGIe9Q+KOOo1hvhaGE
CQagPjXKupFxtnEXcgJvjVHNdMT9hJOBZeuhWzHW2DtJPf0IpxNavthL0wUS2m6w
EDZLvPLyiirSbw3nFdmDNDmCJbEa98rX6xUxdH4Bip70EHSH4qYlDVb68ChBbC0K
sC1DZgFwOxw8wcrzFCzxoouBZyHKCnKbS8w1gL/2zXNcAO00eZbOZtHAPvCO/yA0
cHdCKc7wJa2+OtGaLp6E26ZpSpuK/4KvorpEJsMmnQcdSF5TgzwwLDUQEoyILAkE
cDYqCBLdi1Dch/FNGiti1NjR42dWyEiZ+9u/x5R1nwC6Z8YlH3fHvsLWdc36JJEW
S7uL+jfaqL00Uyb6oqSGlsUyDZxPCWc3rL0LHJAfRwmoedNS2R2HNmoeytWNuIgf
p1T40KpROtYqS59VeP/QcjAZ2EAUTNsMSjcnYiTsQIAQPFKPkGrNjmwVuy4jfoA0
cinWcV8Z6eK0tV1OT8pJgQO+kiwob7kjLRjAXysIykemewM3DwURr8qtcnX6xqsF
I8v6H7WcP0oAikJCunMNGwhkysMITnZe3mxxWTx2EX8zg73dMsMUbcQlWSHpwNoT
4zB/bPgiE9WWe1U/5EqabVE1WEHbhpmhMygVbKCgvtYy9xEY8HidGpFG3OMOukU2
BKZq1EuYHC2Yb4GOTHQAI5rdw2kt9x1nHmpRvVSQ4ysmWLR5zRnbEmiXrV24sInC
WKIQpNvwc52obmPUsaQONMo0oCMIP4Dlc68OQ7BrjHayGYEbsONP5wra7HliTrXi
2+q2E6bsH1miQ0BrXHWmJ/vVdWLBfmWBWCraBoKPb97yBqIiGqa/MF7d6J47SLPf
39gMC7TQKYmZspSnhN1q6s7F1Fw4NTBMvGIniX6lajolw7JiZOpWv4Ntqe4vFpvG
XJ4owHor4kbzRtRsxkJ3SoQecHL7kPfU2wtiulXioYiGQKxiNnCJ44jlgFPlPuLi
ovWGfDSqdWXY2LHL0EB4Rj2U3aIRR7YfaI84cY8u2ZPlRxSlN6cyQPPaouF3aSca
NcXH1kr1PZYgDPud2TYlMjAid+9tjHZBavR/zk1B6BR4XTSHVTkImSUffdOFRULE
L1wQ+AREUq1f3G+weNBMoSJT1QFUU072plAdm+RmPBZM4xCdK2alUj46vaFg6lSH
QaJj5UxXKDB1QUuw7jGOFGQ/V3NVL6EeMjZf+WhLTbWw7gTSnf5cpltOgTJLNQPM
EnBnLr6Zdec95TRsOM2ubTelhWI1gk0oUcR8iK8v/zNdzb+lif7lToECnAj99f5Q
oa6hAf9XdOZRTtDF4XM1yxhMbOyF4hfwn8ngEfvGjO36YTZYCk+4rhvdAvXnMR5Y
QBDMqp1B4Q+x6rxTbilPMX8R52046kgqXy8zMgXXhvRlGyaqEODSuoKdbHRdEKre
fK12IzB3/WzonXIK4eMR4wQuDJ4xVy1Z0NlO8f3LeGW7y2zvRgQf7bEFF3gXhret
fX2GkKAXLJ3Kvz0glnwiA3QcI8a9jk8SY22SxpZBOKUD7tul2BjwTe+Jl+f2Mgmf
Xj5uVzcweuMwBTc9pdRznxYdUiXYpCEwrwNrz20CcVB2CEIwpeFU4frM9eUBjIv+
3uqzJ2wGSkiR8eZZCYzxtxoJnpudoUaPui6WMhEl4QjlWS8pOAM/QEEoGBPkGgxA
SOngtgiPTN32kZ5xbC/USnuMzl3MkxzHuwT/HeTgmWcS/9JraEhDvmaoHOgW5ckp
O5xIL3/x9WnIWd/kIqjz08NwzdiUiq4NNSsMVNIylQSCXfPcZImjL5oZ5lvnla48
E4OMxfS8U0aaGlTdulC0Nfo2dUjx+E6cPkrbto/oQ5FC6rX4HmIdskIxd+yEMvb7
Pji0pnWaUCtxRMurhwopV7p0+Tde5Iy/KKpf8+XeG8HEAZMi5zkxQFg2AA5tgHYh
pHxoyaKBtJ7VtCl01+dheh9n+RF4PbGrcxjF9Mn2A5Skuw6fMgKrOULpKmLZZul2
gcCmDqj57QfgiVo0uX++rjZ+aI9z8GJEEX/AJoti4RLN6c2oFTOCuKP4hFUGc/rE
0jVy2dxq5ZV8LiGRQ5KXebZpL1dFwIk4xmMPGb7yTzisstjctMviDC9F8MhrO4FF
wWHXL64T40pmM/FeADj9/buDRISy2MPU7Vew4JyY7RUFNkCkqFdIoIWe8zepg25y
iY5uIsUXVZqDUvbDXXR1DlZ5ifVlTKQNZWlCikn8sQBp1wSTJsXFLw7Bq9RG/VqW
21t4Xhcp+0cyncQSL3/y2cYhg4qZi9pH4aC+qoLnbeapl454I9scBXTKZyim3Arq
qSiPLhT/BGC5i5Nem/uY5QWhN7Y7C4huclRV9jX2875yO39g7TcBmNh1sYryob+F
zMjhm695R8nnfk2CCiKBh/6mCiTe06h+dbGfv+Gfk8bPjz+UXDirnm6PaEne1KJ5
PC3dm0sMFKRvp0311FFiPZzrB7F0buTkhDISUtTCfLgea75XK+GAQMG+Yb5AxRYA
IgIqL0omBINfsSsCFPAIWL0vAO7cCUGeEObPYI08RxurvKOd753Fg+QPqGzCM4XA
pcwT4pF1mg9e0YTtE0iRek0ylfJQiCzFtuq4zfqG3pdWVvcQwpz+b/y+qQsOfCaD
fqlVA8nq68MbiK5vilsjiqHNdID8L6Z1TtnVa8I7iDLUgPuzh6/amWVKJT3cR08i
JoqNYxSQwC0q3rM1ttFMuFfBNkgDOMkFU70mDEtcPerJSPWXRxWIjs4mfApZzR2f
1ZKUE/KWtcaAWbQ4AxCfkesY4UnoH8hKKZZwhGD+zas9Q32Jb5dNoMxwBCHVyAI2
lLzmjFWJsw81qsNgl5TNxfiJ6SXSkKiC09Y5fQBUmQjx09YNnxLlA1+X+uVGULej
a2uDrT8f+u1TOmxBwm18nWZu9yl6TVU8UEMt4CXEruQJ6Kd9dKQ9R6U9u1FBjOo0
8YS+95QVuDbFJx6V42EpWzOMTgHlpu+GDFFl70B5oukgh4MGfS/goM+CLQFDZTMh
YrNxA8jjmkDwCuQlXdg++YmOw4yIb4ffBji4CA7yCZrM7DMMBbjuIRtU0Z9lAUKm
gipyaBDxsnGEleXUEu6s5XGLplW+zoTdHL/QXGL7YORGQONgG8vnvKS7K1MD7sJa
oJVHdv5r7HWqLMKLPmAcpbfJ0GBPay9JjdbpChzpJYBj4DG+yhA/ftZZwb4WddcY
SQxRBxp+abk5UtQH9iBLBM3dTn7EVHjzQycYR/PLHHYFI8yZkZlq5OYRBcLqft9+
8z5eu5vAz8tCA88V911YVdP+FTIhPNzcnx1m0tHLtPQqz8kvIrp5+8HuKtbqn7Pj
ipnzxfNCfUSo4hxMahHXBViPq9bIq0Bp9aoRaFyFZn86LVQWuzlgkrRj/UqGrqgf
co703Tx28cHUzF3aiihDU7WL7RZ8xat/Ox0LogcDW0L8V12/T3T0bTKjO2KXEPo8
pYQ0wQWIYPgPySugZgSvXyagCRiLtm71rwUEZ8IfTyjwSf6J8nUQhEkSaKuRX+BW
3e1VkdNR+JU31LH8ay85nbt4YnRdheJZ6mxYW5/yVtrOHHhvTCrua37vZo5yT+Ny
YkuwbCKr2PigMYwKyq/wTLIDqPsdochQfAHDvzM62u5dxTO66Oh1NGVp9YvVhpoR
DwD3S0tt2Ktkrc1VQ1E2HrOaHmfYO2jI6utXtE5P7Ezo6/Q5AfzRarnfs2tQKaLk
qpLw5sIjEFvTmw3SGC27nYvnAgY7IfnZjYvTxqtGWRvCj92qsisJrsIK0FSAg1Vl
BzPj42n6oR45//OcdMywzRkIIQ58F/t62B+169ITEAYin4dxn7fEgMbGwy4ra4YA
inIKz5VcCV8+3M5+aj0WYbd0/9m5782eujjpHvUQLadTwT39avhjZbA2G+wa60dF
AvnbBoOPVNnpscRH70ARa7uiUlpJNTJYCCEjfseJzhlmmcN5fX6jlJcophI5E7HG
qpomnra+lnDUOmFBjx4QGTnAh/pEBHZUyq7O8LSQB6Dax6G+7HqNNVBIAo7oXyoO
SjopnCRMyoTi8PKnYi3vyjcH5kdoJDk3P5Zd6DkWNBlYevXvGr1QrB6yhLW9Jlau
gsXamCiO+HBW9bY+eZdU7fNdjTfdMuwJ4ahLQYrfRhyu8iB3bOkwSU/sK9KiK8DL
gVNNXiLBCeFVOKTby4I9ZAorfZtqZW24pSU9UGDCDStDO7WBijH6VfoLRpcPbVsE
43hKDTxEjIQcuqkhpt8DKx1VWCoJ03hzBpI0ryUcSp870ZaHspZoQ4xJ1xIpaEYJ
TOJ2ddPGYh/HdXzA7Sm/Wc4XFJYbnfWhL5BiSD74UC9RT/AaaBZqEf5c+HNAth10
m+6AUE2RHuVF0WWo1HolfWuXhuf628sfVCUNBmJnsZ0YzFbYJEk3ZNCxBEEOR5we
nCBi5kYaa5Hpp3nAmaoPCNvPs/8/fHODkXD5KHkVPJBSwtaUuYisd+hFV5orYNW0
BJpHJ/AcnvR4F5TKc4FDiCKIPlj4zCSM6thGdNFTQMsD8D4un/fNIobx4MhJ4Dcw
+HF0gYF6Jwkr++80SqkonxvdL71kAqtHFRXCqRYQlkrytK7psq8uolub0C/FpsVX
zAOsO48M8CsH2eBEa28vuN676ylF/3JAEedA0NghRWDv7e05y73QEHT7R7ER93oJ
F39x55KxUBw8HByX2TZVYXb2sGC6sWEoohOl0W8U4UoR3LgAIouW1+JKIg1XGS1t
7iea6T6cQAcaW4eioHdlo9ASinx80T6F0jyL+CpWgc6Od5iB1gFqEeBVO5HVitRl
5ntMZchoabGWIpV0qeOIHeXjnt/ciGcEOl+yFjf/cIUTcK9uH2rz0ErXU8bDqVjg
z1PvA8G25sHfHHqDY0bbMOZc9l7XTGOmT/dFc9ejJ2EFShv58nPoqInHoKsxZ3Q4
ClxCva72EP+4G/MLCPU884y0rNlOW63FmymuRhWSpbU/EZT0STK/orAVDOXKvjHy
5iFPpzMgB2OhGav/aZoWEl/V2ZpEm2A/P92N+XZiStJR5HnJEhHU/y/eKvYIL5Rw
dAmmReSe5ESYmLRfK5WVKSlLOX7G3Yyj9sp1sCfSB5766sakLJFvGIXhe+yq2ogf
3BbLRVixWtutLPAwsWYl6owe9VB8jO9YU8AdykoHTp1/c0Bh6dxarjEE/vTQHZ4J
7alKlup4t6jqe5UXyllsMKWihjXk5leUXPcMG7GeAs2nzCCFeBXtQ5CLo4MJaE/W
H40UqStdZ1XZKp/9vGwJ/soXgaoTnnU1u+QaIlhQLfgnNTQkXbj0DojcoK5wSMqQ
wpKw1cCn02yOhfkHKj4Y6xqf4BdENJh6pegEqdZVLkCluH7f/Dttf0USEEflkF7T
rrhpUe7jXiQHPmQojCc4H0WBoX0J7uHThQKBgh8TO3/mNTQjyTtUA7ASiqPpWdfX
nCuv4/8MwYQYWffc1F8xTvC6IE8PQ1q4miOWsrdJgad9eIrrkOMyBhPVlejixIbe
SKRlDhfFSMGYzE7WzAVCmeZPzNbvvZK04h3oGLwtHpXB15IK+9ctmz6PXRYrvbet
VCtf2amoLeM0hdcO8YG8e+fMPwIEBkri5QQGl1qUMsi8K/RzS6KQckia49Sszj5G
vDDpjuUlgHrU2OQFhveHjJON0S+my5ARme1VoSBiLcX0iXTcCRbaRvZjG+TheOsd
Z+eZajMc/HRD43Y3IwZu2J1nD6o/gxSdhLwyn+Xubz1W/vyFGwrcJUcW8quo3BOh
SC1IN01wxv0WvT3IdtHItZSDAI0D6ndnGKZjk4VBnA/talD/0wFPbhYP0MNG1K6/
wGhCmIW43kowV81mZIL/Cm6aH0GxEy3mTuVVp52ioiLh0L59uts2DIUPIuOXLaD0
4n2zHSf0yLgUXQkyfhd0l9uANEcb29G/3K1Mi3iuWOYcX6DfTW+8Sxhc8lIHGoRg
+EUwyxWkAYIcN0MGbOZHGeeuoo2glApo3bJvGsj2GN7XPpuIrkEfF7lIOtg/b5Jf
hHbOhQobUGBwY6NuyR+olnKXndEORvNEQfifG7/RaOPsPm0vygTUSFbHm2YFoL9i
WZJjZz/992Wtdy6G44/GsaGcpV5SbBX9b8Y94xz3MQyq6ryRGtwMCfqZrmd+2oWK
1IY5OLxPZdk2x+3VY33KRcCuTa6LXEkmGQbT32LbmUMWyAq86PTiYnpKN0QbyEbD
ZklJniMvwQqNZYL3kZHge2KDwhMIFKaT10nm8KYJUhNHalkUAR+rfYoMipkX3Mjr
nQJSKZckvLNddpHOOT4iR0lA9g1ksUoSzfXnskRKpyyqx/jHnB+vhZvAZ4usCaed
T1zLv4udJplbceUg9eg03hoBVGwY8b5i5+K3WncP91I2e70J/rJtlHH9rvzy5BeG
fk3gR/716W8y5pRt5s4bhIseRKVUrj2Ea9/hvD85TCabrSJjz3YUv+cLTsYz6PDp
qAwVrLY6/UCqbo47pMH6TaV+wo/4VB34BoK46im8v36iufHcsB9d1+uYUydm5NRw
qqvF5SPaqrjiscsodkbVApcvxVFidJEwYbxNbdjwJ3eel/8N4nBDFPVTMf3td3HX
0vwU/eETxfFy5jZ1gM4xlyD1o8cRohaZqQspZQIcsmij6tp0QDDM33R8TqQEs5Lj
zY+f8gV6rW+jgc5CFQhXCldtD4kUGPRGjQemcHbanPyBaNC8B2dtaxEHNFKqaoPa
3GcDBPMU4S23syKg0stSFQeyHJlbPzB6Grexqw1FWtqLCXtHUmSO4rambOJzzrzC
VEs86i7XHbeUTfHd9iPgg1exM4dcN6lPs7ZsnaQcXxUSCPfVuesqvbmYMU8YuwoI
dtnl1tx4h4aZitn7LdD0eMMW3Bf1z+nJMYsNEm7JxB0t3q9uk1lR4+lvm2Naq033
FJCWtkSY7ptO/i2Z0OVaOmf1wHzeY/IUrrWOcaf6h/iHGQx59qQIy/jr7yGA6Ikx
sBur7YHnjtPmLmClR9pmLQCzHspARntGhN7CA5jpkUQ/qp4JZSOR1mYdzWeVmRpz
vdrxi0gXwNHCBEZeh5ahmpi7gXErrpBy44o87F20YJGL7OCJqOnsJG5Kns+bA1BT
ATGWQkrM01UENebrk9uC9N8BstMkNoFeFdmYw4pHzLLjFc9tuPHrwYEDFyn5PPGh
EJacYPMdQQh8ZNDB7Ww/cyxrgLYnRrFlLCZ2l92ZycD+EpOK2f6kMjRlf4gr4PBj
rPMK7J1LRxc/Yf9WZDbziinGt2rRzizdHCTNhjV5lEUJDFUDS6SX9u+HNFyan6Hr
uXXPz3b82qq8zvKlCgSbeVMYGCJQEt+dmSWMTyXg+2oQZ+7KqXp5ulATQPWisF/F
lKvUqz3rD2Ifyww1VoDPU7Uw5+/mHeDkRtpj0w6aAGBzy2kcvsFRZe5gCeIllkRP
fD7ObTTf4jT2QbUA4vLvvi61DJmceq7YrZwR3sFvSBRto2tHWK4lvhgEW9FZ3R9Y
mU0WqHUVIGuN81j9CiCjozdXbYfn1tyQxWalH+9iSX7noBO4dHnxleNh+TClqB6o
mIdbXeWTHgQN/1W40y1mSKOndYrPANyzXmX1IUbxEpfkxrNZfDC3C/G1zngr2WRe
lqx7OKqvaJHvpHMyJO3q9OXqKJItT4AyGHYxs3BjscQ4WuBEfSTRDMZkVhydJK9D
f/nvdw9BqgOXGOf5nqo1udi4JvPRMymEsYpE4EFXmUaRC5Cnx4W0faY1Ed9FMzla
t4tMrWoF9QMm03FdMEnWKA3i/hFZQrzWOvAfBC16G+cMzRUfS8YEfG/NCfv+hYjs
e7pfQveCLpcUDIa5ZmaPDWRfiSwZw/oqCuTFDefl/G/+HlRozkcdlmipEWcQ//7l
WUpYcqdakcuCJrnP3lFex6PUI6WywoQJMXW3GysO4KlUBr6T9CMIBi7OSVUaBMtV
R9ZStFbwKc0jKd9J8Qo+0hGBEwkcsilugpFBQdPNlg36tNEtJYuBf1i2MkhLYIv1
3BgSRVNFQ4AlJPd+wb4qdPJlTB+ZLXi2puvZkCOcbohiFppQovt46n0L8OFs9eqH
7l8fDbqsXd+gG9WkF+Wae/chomXdixZmSsPmdNCmcZkq1OwSuby8vJTcDBmtNMOD
K1xl29itowE3dw2SLjpr6pr0LyNSLeFRrD4KmUT4Gv/CpZIMwBaWeJUaJ6ApTJDW
nSgdPdpqxlT3MD55h1mcw/1AR/1acf6sh4bJsAZYO84ReArBSbI23vXkOZEgjcBL
zf2ANzNIPDJjI1gD9jY5FXux/qXwjnPSN6VfZycbo786drxEZIYz7VasOtpSIFia
ht5uFG4d50f83z3z2+AylErHUyDjJsw0WtpPBcQEqYss5kZoNPEb50hdjOZ03C41
I6Q/gafvMqJJCsWjAnwW9ZdddVpyqQEsXRwC0ztExchzid649VIjz3d6ghOwBqN6
LgI6r1qebdSCKah4PmaxP+QAS9YtD/VIXhEkrkJZjlsI66pyWQXDLuokzYFnYGJe
F6dGTfnP9YUPIp5YAo9V4ET8KEPE5dy2F5zdnyqSxotxa/9djC0JOtoTQVeITRp0
zROYyje5IJO7YnId+nTpXkLDQ6/yU1yoRndRAEQPckvHWKZFaW5N0OeQIf9Rh6Y8
wk3Wloko3VRaKtzq10+hcZfkBr8LVlB/246BlpWGPRkDBftSpCQPrfgFPxFSkvrp
ZwUpsU7VaGLEIc24Wc+y1Q2gQJUa5JcqQmxr43nVyxXeYqfLt03SzcyXrlLPVbUW
PS/qPDAYnSIJj2xVzlLmuCrmu1J0sx9eshkinho0im5XGesh7sSzCAeeJ9Ze80GL
zT8EUHeByO9V1hb5clt2xNw7ju2gWkV3cp8p6OQSjaW4slnY6JqfLcEbntySJuwG
42wgCgBiyht1jcABhsggkaD+YZjzMbe2oKRMqp2IGHBhQJ5pCfyyJ0kN4bauS3gj
1PrgUuf3hu7ND6lyi+ZIWWoAlBbsIm+MUM+ngSfZbpPAQHBWvXFlK8QenYc2vBfW
OBFvvVusfy7xDjTA7rJ7xqftSJG5zEL3oBrSecdDSOkxL3UQyCYYbB6jpQ7ZUHWy
vzSW89LxZ1MbfT/zsLbruQYqVBTbktLL/+FBmCs4oy6i4V6xpYQn6+g/Z9AmfJxa
671Z8z2nBcUiXEUwwlevrLgbHr5EDyrFrUx0FES+ns7zWVCw1QxzzoQJ3x33CEPy
D+CPd1M/bAbetsR0hFSzM/nUeVFigSs/ouKsAYvjdEAFyFunXIVeIWKgE4hZ3wdR
r4cLQKajRlDLJRMsub4mf2Ilozb29kuOzO8CT/JACzRf+OAwJ9DzPbW8bb/QbuF5
Qa+X1saVofJiEB1YNRQiE73K/6HZDHbp+JEC8rCLMkuBo8WpUYKJqljCcoEC+jW1
3BNXVpXdSlAxuPULxHndo7SLKijfc4/KrpG7l5sZmgsuJu7th5eCnN8k7icStBOH
DPvJo6MjvMdttOOG/DjloxtonQA9isY458WUwFZ9d/GJTvnrl96cQHAHLvENxET1
ihlyq0/yQZ4fjUBSBrxw01IFDEBRMiTIbpvOKZieAD4zxieUkB9TUghRXZWx2DAS
oIR1OGPPZV/Lm84Oa4b6BwOZ+IrSYC2Rl9UwwpNwJsDQl0vEL8EnoyCCaUEh3n1U
viVATpjARWP4Wc3hlSB6zQTWxDuuVVKKi+sqB2PCeR22MFXcb5ISnLJ6Ejt5w4mg
AQ9rdPIv/iyqCJm/sNBgjIvZubbxR5yty6HvlskVMEEDAIygxvQRIi4UShcR8NTk
ixscHfOdLHAt82ahu/DNFJENa2sgrTvXqFBI1+yzkOhEnfSDZeeHTyyzBwlVkASR
NOqgbFhszNWt5PtnCMf24K37PF9MshkCBz+2099FT6n5j/gwrO8vMvNIWcckXYut
U3gxzC0ZJECXlsD5t7ydvl5KmKMQjJ1Sp4K5p8JplWMO/t0u6bu82SC2EEbmcAi9
+zMg9IpTG5BOURlOw2LEoj5sVZk7qRucJftPv/gcB/YDrJ7CwscNw5Bv+K3LulGz
3+7R2JYnchxaSJXObu/oTMMsE0yLBQOy4EH7D2XH8ZokwEE//wKztspxV2aJebaC
/h5xU3ux/04yy7fvRqcHbHBjoajMkgoVyexdAyD5VSAiPVNi31SaVceAOImOiCJP
JRKBJ4Ql+Z+hX47vMDzEmptquasRQiJ9CBnMN2tFkEucSxrfmo5pl1zu2tjBtJmp
AClgHY41S7sHoU5NT2cfFPG+S4JIgpK21ud3xty9ipxvKpXjCylqw6uOhsVfhAxw
UDMU54ju7zkIaKsgrVBK4kcd5b+OQse7aIwIiHeJh8OLeKqk7NXQhD4wBjhzDKOR
6Eq2hryuDKJ8nEuYU8lQxUERAKeNWrKwfdAKdJLaZWnimt4h+XUt9y82qRW4gtW/
anZ9FhXdgKd2omMeHfTtfr/8doWo2L1pME/hSsU+kOfPjpHH4e5rMKPH+i3KAQjg
2YHVOzo3cLukZRrZ6e0Eknw0bnJd9BjFJ4gxLXcw4fiRP1VfZCzQwdfd2Wh/+nXM
/uIcX6INwiUC8rHiz1RoH1yoNAMKrzUQNTtydYxcGT9xYGovuCsVjrdlWSzGTmzu
WvQwbMRjxWcecZPIkfT4p+ZIoSVN6xCtH3A68K1fxfoptMFmBJSEg3AGJcjm1P+S
wUXoBocZIiNmM4H+539ZiXbkDK9tOh5nG7EaqXx1G9DHAgnffAzDOdEn5oXJeqPW
Vdk/h2aHYwhvaMvh2AU92bg+Shr8vvEvXMlkt5g+z5zEvwIxfcNunyO5vgcGOdc3
5uQd46N8ebAGzJ67JU2fVMT05umuIneExN3im45sBNDQ+PWupDTsWmChx3PH+reT
sPNh/jgrGcCybmM2gNQZrXiNRroghGCeJtkSXc5oieSuKrqyvbDiw/vGG53To/W4
lB+HcnrSsJr0tkiSxkOrdjqRxUYR6Z75W+fHTKtFd35SvdSaRU5wM0XIa6uZkiXx
xzPr9784PXVYW1cbDWToXnn3pJC5ivTfxuNVAYAWjZC77EikE0tcGqtHYst7fSzB
Le6wUBaUZTAVGu+dABylNmgbRwk9UJTnQvR/Vk/K8sp1bD/EmCOvw23cApa89NO+
2BUuB5s+BQGLz6Oev4pyDdib4Tix4LWdgFjroCW4HMP1CJIzugIf0qdLw6x23LvY
FTjmyQZ/REkGou0q5oC8WJjZ2uswMCuktCSNqC+fDO3ga99R5CsmEJxQOd5ZCRVm
icSpuXHMCnB0C7taFCKnFWuuui2pfWwyIDC230R561399AlmGlFFhwnGEe3iALq1
2WH2qMN9NldieQ+876f1XnAsVfe16s2wg0be3Vum3NnZcEwRVtWoJ7KggkDLuMHa
+/tj2rDTX5Y2VRV5tvpa091FVfUX+tWn2dGWQsz1o6d3yteABnT4G6+tX/Cp/2bI
cIeuwMqwcs8tDKQkyhGDuCjkv07rYazrY+SG0cYL7ChbTZD3MuHs6pHVQw8XF+5o
RubfG1PPI0kckyx1jOJHrQZyulqO1qBPi6Iy6shLCnq2QoqF/SAusPwImVdPglFv
vYdecIM0Xq3KJiKYoD5ZA+W3+HGdrMDDReh8ttrSrJUxK0ktDvPiYeC25K27qKDz
38eYNattlPR6Mes1rg2jiF8XfZFFAKksKb+yoa/hLbw/bU5NBBJPG+glWUQHMm1D
3w7QWYtISVBAap85aJT7dSXs4BByj6tDpza5bxweYstKWyzMdhUvZqHXRj+GI2aZ
aiG302L5//zxPFxFr64dS2AZjlfUTEkByQ3GHrQDSJg5vo79NkaVEw239s1Zp9aZ
Cc2FBL+SKKgqfWPxiJPlW3uO1BRXPh/dOlnKkA8vFrTAmuCuDE/9IVIXF15e1j8M
TwqLQrxA7Zfz/unYYrR1pdnV6qahyf3fHZ627FbxKE1Y55oLk+hhCAvYgeoEHCtJ
pW5yjS3ZGK0AiRuo21Ss4ne3LTqgAr8VQO3dD10E3IZmo6H0eDps5d3p6YFTqsE5
MygoaS8t1FOsSxy7krNYgmHozdB5a6xPsaMIhbemfBRmKZ45Wr5RkD83/Pzs2b1T
i5OkVNCUV5ulo8NOxQEQG/VJdKgsn8TC1dTeR/Mn/PJ9PRS2HCHX22um7K9qzlZI
4wKly8zUPPc+D/g2g8+voMTWHGeTnimqNlZzLlLNDErJSjvSg+BFxDIg2BZeFHDM
wI5K74ZY1LMJvScg3bEyQ4npv59T1C6glOPQSpojmtV2lsHiPkAbOJKS+iQJSVcn
xLO3cqITQ7bdPq+IpaY3utmdW14mfgUBO9kpqH2Q1zU+Ff1HLHbjQC4NNKawXuAC
q7S+0R817HiP7vRlJGJKdnW956Liu0q66W6iuSHQGpd0teSkITTXhhnW7Q+GsfJv
edhMoiFTro127dru0MtFqr5ZWDmcWoCsK8T5BKQpDbCuGdso2f3dmnUM6RUJK69c
PG5M83Ws7FjsxaNenEuy6NdbVMlpUmpOsZWwoEPlUhqIj8m0qJrZzytkNniUcvm/
4mdCZDG7i9faJ5xIzLnAYLU2GRGrwTEXAZ2Ielj/DHSHugta248JD2EbBbiKmCHg
T7hwWVmeBn29L46EApbgqAANpScia51YpEpYwkjcSGBnWPjthYayZs/8d8Vq1+84
IMJoYyfFhmMnN3dFu5EOo39II4MPZGuc6JWSHkMXgvbqExArSG+y7vKtixfN4q8O
uTk/+tgydri/y+e9hLS1iclhmKAeFMYt5KyplXMxM62Bs2lhr4ly4ulxxOINty/q
kSSeirQP/2yuGF3QKs0rbuAG1ZWgIq6CYdVG6Im18h+iBlQ2qP0S9I+FpePLh57I
/HQibOrZZtwN9MXjL5sqW7ukYsbnSuVGgR2R6EOSyvkrOyrGhpUZMwPK9hAqQRQT
HK85JDkjw0tOrqgugMtbWxlS8oZekM5O4FkU0iYOvTCdQBIUEU2IOBrqmLxZGklw
eS9J3calzT8kqdfgXuh3uvUsB4npLYAREM8wk65n2i9lP3LCiAYIUeixjy047s/c
N/NPp7zQF0huTtjsIyHH+gZwrzw2dvEtNBVJwBuOmw9BMmuIz6FRm7zo6/4WLmJT
39qblYmEHcip4mUFL3Yyzc/xGtAW+UMYyhjfyq0Jq3v9hnugQnqCsWnuiuOnwzH2
89FZ12w14gLeRGG8t0Oo2A4gpFifyyNHvU7WDZxKDD2AyzR6YGSjJYqX2krhyl3P
Zgjllf9p5d2nc2YWsMnzUoyVmjzZm2tjAGxesImf/ZNeGPRy7+FrgyVvA3XWo5nH
jI7se/5RfseVYE08DTBhgU++RwKcuTr4GOeSsH2OppUAsksufiQToGeYcplgZEYM
JhI0A8nDWAFfpIMD+OjD+S6k+aZofNXiQrhmvLlIR87xTx/DlqTj4wFRq6jc3lue
JDCnP8IuIFfARzpmSWXo9yknKxrbbYZ9w5aR4Xt0KFvpE3Qdg59v1hZ/AarXfbKP
oTGIsqEkoorFIE4J9CdlnIMqsagAEBAYB/bMpgAg2kIteAEiQ844WToG0UOqgncF
n0IE1hnz1RQKTO7CU5F+7ohhOuw/tlkKDb2MzTVZgOilFZrjqYIs/sPjP6DuGQZu
ZI4k5kvcc1QebNEbgUN1q22oRHf8b4OXQKVs4hKRo1LQwzt0Ntg9QlofmFqeABxM
hssLlcdyvXtShjHuQNO8LF31c898sp3vdgYYfroAewy/RYcL2eBReEkcX3hwDnkM
PmpoFeagEomVYOj2fQm40fKo+8h1tY+PJGULhEn82LApD9P9rmYLTTWR5HY9qq7R
yxh1UWWFI3ZCSHrGCKHGrIADFd4Y4sWo8L91cWQT2aGz6ECP6eyPjPAGXRfv/lL3
2SyoOsSVQ+PA7QUPhaQPXR/8+hqL6DMzRqA+JGt0MWVaq03IuElH861oF0sPrYlJ
PoWpEzxQWhdMROyQ3sn+7DoUwQpnOvMG4NfBDymbZhuYmGBCjPwmkldYgmv2YFHI
2wvkvjzWlwB4IIK492I92GNTKZKaqwqQdmI4aMv8QshRDenXHINepMmRkPivuDbd
Rwig/6UF61IIxM0rE3QcL/a0QLXSeCJpvhABnejtPYMLcEnm36pH+qj2N+COodII
drALc3sxpkcD2MmvxQN793ePny2fWJUfve7yT0VrgvZuZl18zKzcFtNfR77CyHJK
kJzQ7BvPBPQQqIqtvzh5wMZ4TG9lVIPKfdf665seqwb6jdTpu2QPjM0QfPIT6B2F
xte+3EByeZ0vQoHhXAKoDk2b0iG2lGApWXb5/KdKe4gg9JTmoIcfpaR1VGkiIzUs
5/rOdfNEDlSe2BLnA8Rl8X2zIld45e9462XxLnB14i/0Bgh1dnbJB1CusQJC2iAv
eHRphyCR99Noy1uYQs231TfbUlYVqUEwKlTK4XW/HJZk2mSC6vsK4F+NjLW+jVQ0
h4FK9ZF+ypSdXw5Xfck7AN6AMsbHXCMVYrOM2Qz/YT2Wup6UuWVONNavQDbi/cBd
ec7Ri2ECS7vhgd/+hJ4SeAytMu+5KgIEhdXYzltF1WC/srvO/7M83pbjeZjjta4p
IfzVJCFSLa+WKk7KMEoG9QnAS+1yeleoPmgd6aMo692Is2SanJP/nR+lfEpplIJz
aYzZdHfbt9jSrJWA1HXIauMe2KeuKfcSYp4Q+38RGhVvWS9bCzQvsGarvjc02xcN
gKKDi3JzVampl9a16Cr9R+cbrtQVouJbd1DTrnrbuSGOiuA1qksq5vB2XbydNaEw
k/fTp12gheFGPhcgCiapHQ1MGtoMEIo5bw/EQDGSWJXwudp+525/5m8In+7IuTu2
7cRFHt99LXH40T2b7ULk4tH6qSNG41a2Vz3Va0mU2MLCzLjI1BAKLFM3HnZ0yO/4
FrPkUlnGLbEWGm3bJ6uibUtPm6eWAUioSaEUczslo4tPyo/03BpTrmzBmr8ESHJS
KZ9tnPwBVtYya0i9ObMVzHpxxctsQPdz8uVJlTThuRExX0JwXGRIOTXKAQ/1+RTo
981zZ76LnPdaex0QWI4tR8VVZflUYgLII1Y2TXMzcPGi6H7UrBcNJUNfI/4UXRDQ
YJzkweGkXuxy+JoMekrbQQS60ybYT2IbJhzPcfDiPx8a8f9z7cvJLktzQ8fofug+
m+F7dxFayDzdIpBE/w4NIYTeTqwCebjR53UjS6zedIW/jqY1LARzfkgtcCgH0gk2
e+wDYddapiBH/av1pGcjwrJPvpliDCZ6h+XOcjeHdlkBtTO5ajqLWkgQ/xJ4A1RN
s3sO6yuQcCO35k6FyGUTcs5eh2lWTQrQcicvNGL405M/09dXpHN4zRaGVUokbLTW
BLI8Z4QKOi8DGc70iI+wX46UZ1R7P7gaqV9+zI2QolO3Oma0Tce9wHFsA9np3jVG
lxT5i2sbYw4QXsI6F4RvSZEKRRtoTK6EaUGsMyQoX609r64HxP8Izv5G9pZBAnrE
9o3Pgwtt0JsziBW7PoXcU+kpmeFYfQztTD4+lQN0F7YXvsRcC71Sui8ALhUNnjzK
R9JDhluluHWN3QttxsFUl3Kwv5qgwD2t9Bd507QUfYPApJ/R1Zbxz9BzFXKQaP8t
KFBGOLipXyVR2tprfHrN3FypTBpF7GVX0AXpcYYPD57v8JBvT4WgUco/QKzpRBei
okoTesCyKdRLL1rmM0WEzwD0fJO6melMgsi4XplBsIQFMbplh/2skprzF4yWKEZs
zgyddk+kF5voGovNAMVxf4WuHrsNzg2uQqZAuU/VSWG7YSqH1DF6mvC5d6lMIojJ
rvQauGsuLsnZe4ew0vB1A/lhFs5EydW8ehaITOrByeypqUDrx0EPUWJut6k+IgxH
/Di+u9FbhtBw5D7RzaxjEt/Bc0axrYE7KU3tiXRXTqW5IB2Wu91+U2F9kYLo0oYW
eeDrbaYP1sFo/XwmmPr0woaRtAeOQjp00pxHqPKORLfC24WQcU+ox4jLg4wdgdod
QRN6/HN2PxMagf5YymW6QLjeZ1arqUAkCkzlpx01bOR0gf7XGq79jMrryMmZaTAR
fboKr1TMO4L06VJiEjvOpBXrbPON7ggcqm8vtrZdEAFeEgtMEcpfohxwxDgMbUx0
i/o3XMHSutJjdfOC/byWHGwdLy+FV/G0qiTWJhFL+sU6V5zlnqqC+52uwVvf4085
VMR1YXe3A+I/K725BrqV5O1cerWpPI/wmWj/cfYHy+azCpY4pWV0lBKcyS69/1m0
xn02+dxgAbIXjf5GOp/p5pNzMnQoD0tcI8WIj0hAxFPRgor5o3vOEcBi1DgLUsBk
zP6dKFXR1AlKBqefrDnD83pWgpCvLWRRECwCTtH2a5sye3em650AfpyzXE3i/i7m
+CggUm4TaB4h3CIX6ol/gahk0RQUSKsBs1uLLb/nC1Zu2nz4fCtch1WeMOrW5Lqn
CBoQtgPrX49iZzDZG16wLvMu8LkbNIfUkINCP1nmPlrQYfP9F38S/kD7uCqwqm9o
Cv9NVdLgaKgZetHx1zSf/2HW8fzVfNygVcjrtD0X8p8DNtBrbeXQsmjmzx5xuSRR
lvdxCT3ZE15JQPfOzq0qmQv6XMfaFI8JlVupgvSZzZa8OUVKxZz+X9EB7Y7tUxTS
xOWY7rtx8koFA+80oh58p3gWRx+zVei4CIv5Mc7K/M/Fts4CGDZzk3rGoEvWX8a3
HjUwM8y5v7BwcGwSiIg+J3wD5INen6Uc08Sm/Tm0JaOK2S5cVkxWxtApvEYZLXL8
/ofhfPkag63LYNfO/fTt13p0pLOd+bm/iV0f/cZX/VWC5d46X4aHOuZGpsLy3qds
CfdjP9N8r2KeRDPShEXUH3maH+Q6/RyMqc8VJZ0h2TrrSAom8XDqdpFruEIH+NRg
ID5w6a4wwvtPxrdKSPbLpJLGYokEHzs8RLelM3Ex9o79j49rfr1Zb1xH1JCO0UYC
OH6fKpRHZqy+aopkLS14q0e7lirF/thyzmKRXm5hE7R2bT0mkDG0cMITS0ZMpx0Z
OxuaXBok/oSV4Qri+3wPJQ8Y7heBJjcVGCMNBrgsm1vIU3EFXsGMS/wqY5bEloif
tRZvpUOIRYrij6HiIdGjVY9Gkz1xeaM38yJosPQciNDyRtjk2GeDXKo72nrHr5jQ
svgLxxIreN9r8Z6+GYGHA88UPVstfhIGNGoBETUThrR1T2ORmIGpekYg1KDrubuN
yvwnvUFWE4+6e3wUhjwebPIb4xYh+5bVDlP2YzY2hcYQ/Mf0Y0DDjgUpA7eu4ZTU
JP4lFPfOm/GR7GoquWpnqKMIM0UpSdAQ1oCE4TpsCw5AUUlygS7EZQRRKLPPIhb7
fkDbDtfBnd+jvxC7NJEOCgfMJ9ruuwA3AS2DVvVP4mBIH8/Uh6WRTqs3Wc/h5eZB
jm8/gB2vO5v6aufh+iollWwTlJxkITC7phEd3k5MLEiPr45klvVdfvqip0/gNjAy
KD9ZHz7I0s0SUdTKvvPJzKABe+6OqGLNrgEuWWnPBTfNfllfZ2ZBJJNoI49VVeVT
nmepviEog38osic3TecLXttBtgLgrNYFl5qIkB+pihWOnXDv0TZyz1mvXpnzG0VE
DyCYvQ0/mVviZSxCVYdXh8Bj4T8WEO5QtyUJXse+SRGExPWVPWGqVi5JyPfb1pTg
jRcBUmyEOZzOC0H+5Pon7JB+f+JHBrpjLpoz4Q2Xmjpljk8kP7eICY2xWm+mwPXa
i01LjnhbkNZL4O1OoJTZaaWpvtySWQOUPdeiTKQ9MkPEker7Dm0OUfXBLuAlau7C
7CsH3ccxtihKP0TOQnNJ7x70KJizcBbgzICw+vap06dACCXPlVPnv6rGrHXJRpiB
xStjrPFlJcSrsCz9L/CPjhHISGTJLD6G/wgig02plk+XEDJHChXNmC3vz8ZYJaOj
yzbg81xX/hr/pOhYCRqksGoys8fM7TKFiekABtWnkg+8GjbLjscNkT1rOgxo/zbE
8xBIX37iZvWx6+TC9mPqutaDw+CIDxdBUc8JhmBx55ic/SuJUnUn+hq8cCwhkR7m
h8cv86/qxmixF1WoOskhxDMBrzodz4UQq0R3NMUsDv7CF3k3/7Ta6tx8cxtxpn01
hj5H9B8IQ3ob+ZSRWV4sLqtXS6Z9XWpW/FHN9SgZhfsSkY+7F9N4PtuUvWiM77x6
jx8oNzXjQ/rIROJIW959cDdCgEMGrn/iKilgRomMhz18C/P8q6c2nAOuGGMBAyaa
mI+0FbDV229P+07nezXocPp4QRSILbctHxK8n79fVm3IROLFotdw8t2mSMRa8uah
CRVi2roFM8nCA4nzA5hGyhcaOZEQ//uaQHnfvb2tPqiK7EtZByTEXBPzzAbooHwH
gNG+K/bI6fcim2tNQz/3UVL3Awy15fvRcV4AgDOdB0iH146WsEcjshEK2BIRDdwq
7jreVI1/5INfiw1Ci7Jz4ZCyda39udJfV6qhIQ6Jr83fM9q8LJyei6wri7Qf8Mf+
BFWo1ZWkKsPmDS1n0qoqIoYU1sfl2GPNX05cO2gw/x3HMbrK9d97+YUbiZRVqe9O
3A2GK0nKAOrETlI0u1IjdLPQFtgADY84dTZY6V0E0JXSH7KFowJbtkWwFEOB1XIU
0+R788eGS7lqydfj9pH1vFEKWGtff6AxV7+EZu9yIW5wgasTgtJq3l3Ae7jj1LDc
DSkBufvwFhZh2S2xd0xpySohshyTKAZkqXLd2oLoWMGtVO+I3YmVZZGFxx8o3oqB
sAn2kP2Fgv+QuvYPDjD1qDQB6LJdgfRv9QuGOfb8oMsefogoP9mA9QZB8RoxBSTv
sQ+Je5HcUqeTB7uYy8z0fwvEvVcpUh5hQSA3lmC/MRgGNrT8Ti7pM4MU0JlnjMQN
PjLEaBKUV2cmObJBbdBf/yUUmQUfbdGuhn/xlO0bd7wn087c+RecRlVznjMH75nd
Nv8ob50NOMo78ztWiOToCLaLxkQvXw0rZy1qfW/gcswmdkVsoEJjetCidloAYcsm
VtPFuwOVgNJnEhdkEoB+LGPvssk2V/pp9UDuuTmNwNcM18RtlbX7+VYwrLDAnKB6
m7D65fnzuzI9S9w5k7Idc2RM3QXymaVsGOq8qfnzXpPAIJLMyqEQshIn795KVjRk
Ry3Qwi2qbDMpPaOhu14tjFbbbPReClR6EdiAv3X+6z0YuaeTmmOvZ40C904IkMK6
R7nPkF107fizU4Ten+tPmtMoKypO7gvTszNen9gx+pYwbMuvs7JtWjk32/uWpugi
xBD17JOQlAMNv7b3b33hklZNNUdDvHvijpzVE8t/osaV3ipl4GBudkfo96MTHRCP
iBpFwxsrLcm3W85pRfVITjTEQhd3pSLQ/blosB1IKyL00IPELxfBtcaUJ2VNAOrD
DwpsLMqUAQ55ioDrSw68M+iX8zYXpiHiZt+1pD/V13tYSZjidF2oSO7I5tSmkcKJ
oGyz4xTjglynGelGGQdNjDe5p9/ktihtlcn+eQPoe0r11ZCtjdiGgtn5TkqF+GY/
WINaImhUgALFPuc24RyjTcoiPJg0avBO7F6wQDIzMz8ld3Xu1bGJMHMoOI76K0Jm
/hsuaX5dZnywf8OCZl/XXn8g5mTmj1SouJam3RfSCj3VjbdPRkArfofK/JeP5HgK
14Nb3fRrkCJellZvpxyCgVRqXlr6zPUMnyxp6kBJlWqEmRfWMkcXBYrWYgc2QH3A
gaZyjecOdYyHBVvfuvwB87sJrAT3N97JeyTPaIOfsZStCODgd53xSM/edxwkwBMc
jvVHUkGF6c+xam9p02AnmWfNIInTrGTdDNhrx1B2JW56O6GZVs1bVUAXCAAh/2ZC
Pl1jCYGtA+QM9sbTvkxpzq0kr4c4lEQhiyPLZzL1D0CdL+IfEPIGowMgrzp3zP0I
BOTxTqZd6mG87H6mD7sbWN84IiADW4HXSg37yzRm6A/tSIJ0GiH//ZKVf0Bs5E3V
Kq/UtwrAYKZeRKiEgMOoeGetpg0siY7gHlrC5Sc+A0GeSdZZRTSUXNfhBT+fjAui
E41t0IJr6E3JFiL5c9fr7rElraHQDT388bLWMwe93Az19ZoAzF0JCxxIRh0haZlY
4tQNKzbnMMui82UBXjIYoUyu8qj2z+WtmZGwP1ro5/NpdPoPDIua4FL/A/fK6k1m
UCqIDtVOpa4ZnJMipArQzGAdtVlsLW9Dc1Mk18WBm24fx9THEITNFskYuY1eWJA1
bnkXB+/0XM8MbUvkPMhkKQCdU+/ku9mVt4+CEWOgjevPfU+MYDpmhVGXHsaLl6T6
Ciib7iQSby6yWiTsU7aLaqi+UDe6lLU1jAZqSPw4fuavguZzi7mauY8TglLxofWO
U5M54FALDRdTm94rRCnw/Y1oNFA0DwUS+uOv71tNwScBYm7zYD8f5ZCidKxhpqMn
WwJgwDYyvh5azcu66wsfAlGL4IkTITniaX+aH+fwJ6TyVCj6RsCIZLdcyM2LRPPq
88IE5gZG5kuBSP30nAr4v9Zh3uwCtVsUmKBrYjEe7phVf7Gtl/0WVNjaTjIEMGer
tPECTDaKCleM78jeWhr6uG6bPu4ksVP0uX4CZ78WAWJaEr1DD2bOLy1o0Qp4BFnt
TaH+UxE0hcYQca0uYoDDtfomNadnDLqtRoPx9pijVd0i/MHauRwTvOjxW1MGnEIQ
8NMRl+xRC49X5jidnMiYhAmMW0EAjkKoywKEs+/MFINRn89yOZKApWn2ec8O7M6E
8kGgMv5sTPrK0u+wQNSovZ79Gw8idAclSaPFpmEkut/OBp3A7YkZpneAQnfVDvKF
DP66W5Rvb09EEI82XShuKehd06jIOHbAvCAi4gvscLNFUF/QZJEEJV64zAQdl4Ha
CQCOSwEGaxV0tIgC8P/6PUu6caC3rwawv9o56nk3C+PnjS1DCRHwIotRjF1+cSvb
MjcygfgSLK40w2TmPMIEnughTjhLkDEGgQBWfJdHwPk8dK1WEOnm62Gcxban0vJQ
C+3lNZ4qnABF44HhJW647NxnX+cQofl9j1PtStIpWfZ37FfuW/rx5uNwhtL9VZUg
EVu53oHQlmgvFTjtOw0xC6OSWTc8hn+QGnJLRv1SqPhoN3XzL89/BiFFS4Es9nJw
tDVlkXB5bJ/ndotdmMOkRlbXHky+Fs+TIZKEUoQsJzXqYXuyO2q6CPGoCu2jCOlC
mwSt2v4EAmxSeghL6G3UFWIjnVh5oK2/DMvVGj5sreUBnUUAQIrbQUsXtaJX/8nm
HUVZM+XWptOyQhqsydnFIhapsrNpKtX4gEgcnB4s2ZDPuFL1uw8AtMA/1FVf4rrD
QzrcW6yZIeo9aIR7lzVyE+J1yVSVby/xm89RFrnx5X3Lx/5lX+w40AO5kAoJM1QJ
iQ8PiryY/d4aZF/FjOAaD+PqdqzZK7E7XcZ7M2C1L1nuJXQPB6CnySsPDJOehLGO
glM7/rua3PBYUf9RdYiQviXK0pOz/RMlYIif90G4bSXB+C5GjoNu3n5rEJf6OmNv
dhZ/vdfEip2Aq2UPUKKSx25uH6nZlro5fN8R67A97OS2zI7MMmF4Pyh3cEWChG5Z
ecPfAVF6opIc7ae2LNgy5vh0VspR3i/PY5eu3C1kGFTMG7VDhjtNhCngwmNIzRnz
o5rZ34CDzW6a1aC6FMq4OkT6z/jdaFdD4VmLDvRCipM+QMpzdCi0jhoZOpJ1Z0zl
qmbbxtSLrFE/wnasiAq8BNGhLoamcr4wPDFfv/l49xDCMHzKRwTLcPateU3Q0Ubs
uTG0B2QhYdE+LEsf9HASQSgFpAPdbgueOTabzjR1giEGq+OXmVgQv7dKSDDO50Ft
M3vZmMdOfU/G07WMtqbAKpvop4Hs1lqq0tO8d5qS9V8Gue76qBs3UU5pL35si/AO
WqBFrOHN2mvhHasiESlhheIogirnMdxUmGkJgtfeNLCzR/G3xyy1jCOQ+p9jV5nv
0oO0rUs5QN9lJhyRKVMFy2a8iZ2Kl6eP1SlUxnIk6aNu9VbMP4FawlyswAcfVGJB
nm3sll/PZrEJMu7UsIjFZpNaNnEAcHwUFAEF9EsdCNeHV6pP3MKwc7CE36R6nZyW
OmMO8PDzLFaeFzYrQdRjttm/Dq1FwUVyteyZ3mq0Epcvn3Rc6Wx1Yd2XQw4wmkNZ
bVUzazVoWMARJ/BaKIoITfJx9x8qB5eePfOFJWsnW+9UBEgdIugCow2uFuS1aUTx
K/8nulZA9ZSKG0HL6K9CGChYYiIHNvICSpzOQwqgcXp05rYx3OEfTW00z0OLgTLk
c8ghKjhzic7M4ndWa4YoghvJA9GXx+rqM38g1WL9my1rpSmSoUdjzzbdjvi52yUE
48Il2yLYkxDkS7N75RQPRrvsiRBo8pNFOsK2fKlWixCs+OSxkMmIpi2uq2EZi33d
TFvmovcGkil36jAfAk7iYbd2XOQTtRBBwFClj1XujruUfC17/BwTbZ1Wovzjhm6B
A9hZ77hSFwqScpoBEYsje7w7k0duK+J8WlmVe6NJ2P1AbE8ElV3Q2IMqmP8uTyOj
uZ1Y0CQKEdfNRieJuDo0/WdO91HRTrDQHiHGVzh0RMR6g7F5Um/GHJNAt1KCOXgI
hkrjTe1zdzKOCjm9SVkWvehqqG7x4veFeoY6nr3HlX7vSxAU4E0GkT8U8R2z+LpS
emsJQyKufWf6ETfe3mRVVgWTTRogMDrXXF6T320DVNt5j89IerQKdpwXOII2nClU
FGBEF8y5CPm8JIyc+rPfCs0Ho5t9yO7A6chzNve9Xygv362YNKAmbrQQMil05qhf
pukvDd9qg/bfFvYaazhIqykGPC99CqwudpuU8iJLTcreO/P4WxHDuLlniOQ4M8Lv
qG/ZdZbt9PqgAJsbTPz+4Dy2AKd7XfwDcMdart3O90qe+FAAs480tWi7KMY8BhH+
70kNFpvn1fZFoIHE/zavXFpOPfkOYr0/CX6irNfAMAWOzdxeY6ZMLh6SD/t6r4ov
witHnBmZuvwgRDu7rFcxz9uje3Yk5KwWZKLLRyHvDEOEcjrJ4gQIKwdgRRwF4qi0
nVfKj0hxmlQc8chXYUurUN1lLpvjf4/9huPJ4YyJZf6WcE1mAX/SPo0bVMYC8re0
tXoY98C3wAl61CDsHGGtHemWE9ry75k/rDD8BwLxReupEnbUpTe9aFF/EA8YkRdT
m94wzzO3JkSHVdKmCFAZDl4hIVswAJBzfN+zX+Hsh4Wh6a1QJbYcjUK7oRY8MXSo
zC8Ka281sUDOaUeOoegdyuqeMPdfETv97B9/tAWb2MTlEfhfVhnCjzWWM++UBsZv
/6A1CMLYf1MXlMoWFN9wVggZQfSQXmgygL0K/Jb6YWxTrdlFqP7B/9jhoYzXy5Ar
bPQHZb7lBkAkyrdGSU/DhB5PGfgUezuUcYHYmVRoSIi4Ir9Cmc9SQde261zQH1Ov
cEC2PZqQ0DHNqBEjVxsmuZWHgpMqB3G+/x2Njav8BkiT7q7emDce093pO8+HJX8o
kzRsE5px2Go3/8p88iztdYRcAp41Q4aoqmMJjy6k1ZDd8VtiUK6XanRvPSfwMsPe
QAQWvxb2AsXOo7o3Eb/PrKhAue9hXFvt4B3oMmlyzp6uZEgR4ZzzuhEenirlBEVf
3d/ZGs2goU0YEO6b7b5WCuRFUIPJaVCVxcafMV00KhDDvf3/BEDLffadSA2quEfB
Oz2EEaDTsTut7swqj6nQyoTXuxv/if6bMudZOKLMO6xmrZFtq1cbRSF+PyhqHE3k
U1IjQ5vPxhkeimf1Gr7pgVmdwQgj5C6R1UjHpIujXVTg7VjPkP71EEqOw0jhlKiQ
Ce/F/Vj7yfJPA/hCcsrsTDtQYcHnA0wx3kVvsghdUKUXGOLjhiWEI5QGAN0CzZQX
qL8aW+JF/nwvrtbf+DGppXLt8OeI6Y2XxzkB/tqQIUiVVX19HsUNa0e/ctkb+0E/
INKb1TIlKWcvmsk36hnLr5Qp3iq7Bf6UDQad8EnkT7LcJUuzWmLNY4bwMNF9LZC8
sjLRBZ13T2IqySvKeG1GQjQi7sTg/YwBaHRHvMVAQvh2RRBI/vkpoKqbaCKHUJXL
g8ARsOFeMqtE8h/W+E95OXD1Jc/xHY7d6wz1qxuggmR43JljxiCaOMy4524S2neg
qIB6u3UgyFBHHr+Il6bbcoz10iBiuoyFz6js/av+PA5sHX6aknVfiF3ddrhC5xtG
pUb5J1dZ3OoGjJWiWXq9SamVMGSlVP2ThDyURcnjpuDk+JIFSyxKpa+NeQL/KBNV
OW8yytAUul2xCh3SOGHk0jv3m0C9YozVfhb8/ULFoW5OUIr65z8M41TF70GXN9oJ
GaUEOSDaRk399NyQC7LYiCuhyLu5AlIR3g5qWnevBnmD0GznU9e6Q9IIxMVHKL4v
lVS3WleCrNGON3+ROqjUtUp5dqIsmQ4JvHnjvr0xtih+/WDqq/oe/SVnlhYDHsxy
EyLII6Ad8k2FbTGn4rlyTuaJact/iBJCzkYdPKVbdHfNHoaFXckZt4kCHEHpL8sV
yQPBqShZUCmSsHU6/FEeN02qHTcsAHd+OiJcr+qOfN49Q+VM2vJbr5KuXVSHJkX8
ab/BJinvOmaOmk+A5JpBiJOPbf2rJAyeMuXKY/YuisabW5+I7v1X4Lq5uGCjnffS
3YaKSsuvJKF23QGu8f+GHPwu3vdG1vXxLZheHFCPFw2+rhAur0pedi3dkh8l2/cj
iKk60OJ5/htmr+uTbojNFECKoUNGZMLUBMEiLq6r4K4BvMQMmjEEYBy8yY6BO5jx
FaRkJRkEWonnCz+7ZEhX9pjfmkLcR+TDRBRgpePA6FUN1KvmkP63LmAkcySHhHC1
3mUF3dz0vTU14GOxYFqG+9yvF/jJuT01/Y+U7OqQjgRZ7E+yoOv3yz+zt6V0ct4U
dKgLQFtQ2Lo6QfRjKcZLDBbZdGdiCrvbPZ3tb9RIZ7En1Xt0YICdw0L+Sr9v4bCt
icZ/zRScDSr/pYE6jKSG0FM9iiupsEKNJntr59zn9pe83jMkAX+T0rAK1dsUnqO1
FSY9uSeGE6Xjbjy3BrOOLPrFrZ8iuSy9d4vXWvpLQhtZ/uGX/ZXXr0FenpHg7RaA
RTPnOFIjpka7Yb3aHSAf8NQ89T2cS2jyApUx8wAHCZg+h6RpkRhVAxWU6Pw+2MoM
zZ42bcMrWY4kBvYK7sjjbr7cY2a5dVgLZ11y2fq8gDCxAI7Mbz6aKI63797ar1CV
TRn/JkyZSu/Hra5lROLB1I0eUDcn8N2pCr/8FW/ur7q2pHC2ubHprKcAizXAy7VJ
F6DKqg+bYOyAChxTHkpDS7hMQ1ph2TSNJThHd+qW8L2dD4knl0S4w6F4/r0h6PYh
7d7adx7/G+TDfpjhpiA7BnIKRyKEmGyDA3ggvflXVnklJTQUOwd1isvNUSZlPx8g
CR4ye4ik+PTTRBe9456GwJHkxYLmNHFSds5mMcxrIzQFILP/H42sPPYRijHjgll8
fjsvoAfPd+Ks1/SPIRQXnGc+Z0SjRo0JUpm3CIyyjrS+xJqZYggZuAQkwROsKMOO
o8It4rkIV/9gTUlUPtmbEJCgDXKdvEEWhYMw85++kpA/b9/NmHXin1pwYXsMoEYz
bprqyUXHSlNecOvVyasdBG1UpkqO1D4ANquQNtBpXYRvLiDVzcV6xkWuGr/c4NBP
wDRn8r1E+nzpX3K1Rsa2178rrHQNwNxP2sigLDbPgK7bMwPYTO9D6wlgLyAjxWL9
6FV+NJMU7H1vyqIteoOI7lrDIEblXq6jxFE2VvyU42uC2IptDZI6lU+CTKP7X6fr
QSQYbXXRtUlxRXqKSG07eSTVNH4PL9Ots5syBa+ljGEbM0vF2sH9Pbfop8etzMp+
pb4G+nHprNzWkmDplV1fc+JX8sFbNK9dep8cTKvwmaT1P7me70eiwbV3+xmrkP5d
yylxplyRr7tZ7xOyUp8duUe6FssWutDcQQ1O0VFFv4oKnp1MR5cijoVqhXK46hNg
32f488bA005nX/67Jw8/QPXvHbFl+usAyM6Jm/Xja7kQbgJ0S7xKSKfT5OA9zu9w
D9GGhXHLbQ8tmyWbiNFkSy+pqHHZNhUkYotb9tpJp6NKrOtaN7qE8G6KGyKS2f3F
Jw2VHIYpBOpncS/vgiDkF/72SrmEWX5fersKcby1qfk0OE6kLI1aUFKKHfux8Cxy
G6fFhGIdSMnYI9HkRljnUdwwVTGS7dGLuz8Mu+KoFn/+RlDABFQAE3iLoxTK3aI+
Kit+pk6XUwmweZOVnllXNLvAU7awpFZv3DIf0UhMZkJN5mDFcTZh9IAnDIQGCaMc
hLwkpjsR34PsKlEbJAKcCYbq+GigmECxArjgHo73/6+taiaVsFryvbdpeSMJmGEo
6vg3rmOePx3pxnolDfv746iDfvlCNR8o/0JMFFfKnhjN0vmscvAbkEO0nB7fnEyQ
Vyda1KDB0nsYnOvI94EWpLgX91TjkVHwhVPoKf4RoUTlBOXQXpzOSieDNdJVCGQZ
eMA+qSB9EKiOE38Vax93pyDIT0sA2rSt2Nzy8WtSLeQ52Jtxur3DRgLEzVKWNZDt
zuAwFWU+Mz/VdeoADKavZZFORPG1RdNwsfL7zXtPImlShg/pAL88Xs8yvHGqCJfa
qUjFxK3ARBn/qgCuxxlxo6ltZjL/VSDdtvVuk6M5vN10qMsPTlzx6zYCgTD/bdyV
Zw2QSrDTA/AR6dW36s5sXMS8QXKATNeaV1dld2+I/9Yy4/L1OlxozsMU2ecCZpKH
wHAiKegvm9Kda3oPEae/bOMj2H5lfRztfbt+wit+5zIW+X/wPzve8dHGfnvp4FZI
L0RrJrjWFJmLDc7h3DdfZJ2pUHE3p57bgammv31ZBkIx/3bfLjyB2T63n5e7NqbR
DNM8HO1tr4JtKLp58ASIuCHmAkddQgztxTfjInFol0+5V7houoXxiaBOsfj5nV66
f2J18+2AvX3JU8RMf/XLen+ePK6egcVFWt1UrOUpvFCUF1y1jyWfN7y+slaT7kjs
WbM4S6R5f3B5avrQy2PbdQ9jyWYQP6DQkz3F6FAYogauV7tjoJ58hHYgnoO6Qg4b
MBrh1OcwpCcdG8dT780MjBPdVCD9oviQIbuHWSbpEekAkhI1NmXMYppDrp0P+JMi
CJaG2F5y6ZC9ZNML4x6/x7/qGk3HSmFtfYrUaAPCxXJPD4z3CuvcPZiWZt4qnjyc
fUAZlWEREdnqtP6mEmJ5NfuurNHomnNj6MESqpDX3nRjEfdGEBAaqkWwW4iSVrOe
jPqtp2I1iJ3pqb/PW3qRPUvCRAuY9d/KosZU9QhQ1ElYfhP90e5lRvCsmttw7Tt+
b4zYWXty+VPR+GzNYXpGc1PgwmUpHLSFLrXZJsyj1oZbPCG6T4ejPIN9IwuLAw8d
lSQpTUAPkL12XMbajnaMqzAtoZ19sGKsBW+jecYtrLVB4JARl7P+mv/FV5bnjSZ8
Hhht1dfUp1uVmfZfzK1JtCW3ElN6zCOlU1kJV1jHXeDLxn7A71R0tLpMz8NHFbev
MkESfCQShPlr/GzqkglnlY3YuoQyZYIj5K6gAI2iXAt8hUMxdxkcjOl7XCVp1s5K
vFF4jlPqvLr+ACZ4AyYlB2PVadrjuaPTI9/UxQMWb6pPHV3UtrhgJGMhoH1Tv2E+
8BaTWGIPtUPmoX8KZzR6RMdI21lOCJqADZ3QKAaKUzC7UlGlL7xQS//Vd7tq6pmr
3AFz6hVWEXanmg45b6uyABDYPRUog0ldMwN4vvzNcv2pxdwTKL1B64KKz0/6jqVM
41Q409aPgD/oCTn3eThW29SXTIMaJPGjdd1/6IVsm2PVVkrcQ5uU9J+M95mHmu4x
YgYufZkVCZSqsH6L8tpacIkJuW/ql29GXxS+Q9Mslq385I0j8+VxkeiNdHzfYCNn
SiZzexaQkwXn50YfMtNVGqrMlCHPB10uf70jOr0eKSN8Nk+FHFDlCpeo5bviIgnl
DNunoR6XjYo3ZQQoktDQCBUZcMgP3bzuokTZHnVC9+sqrTER8IyFba45nviWVwfE
FwL9HWJs9Ip19qZAml1EbNQzJpg98R9qKjMRjy1Xaixy1joY0XRu0dmefS8JPVpx
vS6f06MaLxrR68KOWdJScq9tAzWvIhisVYK4KTCptRmkfrPivyYJ6ewhlEAZ+plz
cPdKu2S3lOLpRRR35V4sNHjh7lvX3ForMX5UJnuXvShXrHNsBfVM/RXuiC3GSQp8
wKPhImGBszjv4N6+JiB3qaKsAP27HOKsNSP4x2KmFU5H2dS9FElED06CekTvDFKR
n48UWBFRy4qa4DHOvczOU+s/VJTOJHNYFmapDemxTX1NPfSknf3b9oDR47Ywds47
vpA3zQuIrWR4NuafHfnVn5PWmZM3ZnKl0D9u9a/McErzfYLV4WtH+J8Y+R22WtAm
hJyF9QeUX5BjuVptQDbWGv/ooTfPOxA7eBE8bP19jbaDNFPFbnfSGoCKAMbEWB6d
CimGyB9J0PDhUw2aS2aVoz9rhNlOGUqg4QPUDB7AXHFCl0zi2OLIjFJOG6OYmokn
k916+1DtHn9++K4AeHNvgDLdZotBtiNIc2uZKLZq9eojhKgwhYDniC+2P73tIYvn
Kj9If4uvounSTztR+dz3lxpZso6dVUTlwss+cDC8xRonYW9OOGje5Rr2KDh41pON
Rs9xRrXR3NkXOayLyIzoU05IZNgSZDKnwcYx0TZUuIdqL7f/a8R1Bomhinevpdbd
74vXkzEEwE2gr4oOihB9WQSuvbxggG8ffWgIXIw5RcKQ0+sNgYnFKDg/ZGiwmjW7
CwMUMFOWqbU6E9sCeE66o6YHvInZN1rv2qi3J280eiZkR9yBahu9rVYr/Ov3kDIe
kDUYE9e7DlURimUU3ChYMJCSUMb6oiT00tEVy+035PAUFdkIFK4zjWaPnkAnC7nj
xWWsPT4A1DS1137Bvgw0jbhXNENX4RfKfjpbKBbcJm9waNlniA2ErkBUqBIGmBld
2oU2JHigYU5tI9qCPomwD9ZKX1Pbbt67EBE1LrrzQzVjinmoOptjQUwVIWylf+Cc
+E7X5QEtXh8akpf2UcGq4yoU4IpRekP0VaAXBqtBgJjC3kBuMs9btxkBacS73I/+
1dmWutfaUX/o24ikEat/5WmVsUkdfNDq/VhI2vi4uyn21VPDjY78Jy/rC26SLoC1
87Db7IC+k0f762XbTNQVTZZwlnut3kxS9ZIihcQh0bJyStvSZX8NkDq01H19fEa3
kVAoTzmOheKOG3DLGs5jAWTjj7LRU2BPlNIrhn6B/Px0NEoGPRq0IJh5qMaurIwm
C3kAu+Y0aoDTeLlZ2wpQdMdgmzrZdHZZDny2YCAJSJI53BN9+U8V2vOuFnYPbqeu
IGkJFd4VhUaWx+Oc8AkY8TbDD/hm4YUni6TSXx/agnVcrjdmLlFAYZdFAOIKbAhE
SZmKVNgOCoe/GG4kk4+aWCQJXcZdGezL6npCOO+NGBvlepm6ntOw87xeVyYxUA1P
KF919a0lZaoxZczzKyXEQ7T1IMxXadmLGytbpZlnvlUbeo5iF/V1XoU3LXzu+R9l
Ft0G3VFNNkd4gk5EM8B2LekwpeHSlZ52m3gVKTI+2ZkQ04vLcfIgsUcR4ibjwqR7
0OoX9LvUzhxl0PtKUCffRwysD9NCwQX920gGnN2n4I9EPu55nzzcPxt08965kphq
uopYZzE3SMANbtpm0HduxYVoMzLJz26e3+F7v/Gqpao/x0yIF/SPzcnlssv5DfUO
/DMqvm4npVwvp7qcQV+W3hgrorMV5ERpVlPIyBXcQaA3uXg5d4TceVZN0+fY1JwU
oHerc9hRlYLtS7+U4EdqkXKtny5GYY5Ez0SMn2U5gUqNGRK0D8vpq+WlKv9g+NVu
EWJg3CudnwU7LQOs3cLc1MhsICdZcNmY21qMPM7HVfolCUHGWHaEA1GnxpAVxaLO
oS6GfcR20q6XdlJ9e2Deb5efPoEf7TuaqD3vj9rYTHY4ZEA9NLehgDXwd2gPltl7
bwnoQGkm7sKGw/pK1fPiF11GVQ7emzJXTwJNN1nmrSkY+TETvfZDWdxu77Z1iG/f
Oz96X08w4Ee5ZmgJw4IrEcqq2M1Ygny4DO8+4avbuS0AbGugIJidzyONrjJtMc+G
wX3bUdlhHIUkjpSt709NKUlkfyRuFCY3K9xFkDHnwfAaoxOsYxHjX5NdQBBDfgRX
HwaH8rHuXArbR7rqVIBrXaQq7HGCPdhotW6ZQIU1sia+cvNXQCqFelqfR5Yi9Hol
6xPK/27NXJkIWwwzC/XKQwyfrxOrEGcd0j1TlIWevl2+MX/zGpDRR/AOobxZ4x0t
17klKOlXrHAOFu0b4y1RkdHI44L6lZfOM76zhI9uto3uLfD2RzVO+hb3N5gdb/7+
fEwg+FRtLRAgSu/KPj8YbW5z/sepBtr3MKDVGnT+3hPpfdC3mGOIeEQS2n0MfFS9
d4brqYupMI6dhckLnqLwVrkIYIAb8e4CTVqB4cPI2TmpFogMzmHhivtAl4OOk/L/
xbhd4cX2zyIoCWp9EapndKcStyAxWo5l43LVTsfboDpoZhOr6o1JBnll+pYdtmEY
3jFOqOIRRqpu/2nbsCbKtVAO4fuk2fCcICS8SZqr9qxiYUqwYrygNpyJbv2cLQcm
yk7diS5FOKMd8TmxuzTSgc6d4jffMtTUq0hIucdhouhSgMS1xPCBwaxP7fmpWwYv
1lcRPB2ja+Ie7VLMIJXhFJvsgA+ow+01Bc+HxwXf/MgqBI4Ra1P2iCvoKF4Oa2xQ
rD8Kuc9uKbbKVgpD6Zel6kXr7T5rwDv0Q5jl6bOKcgBIcfkzPy3cqjYzUvPIog4i
YC3RJ02XuEJ6JuqgKrk5e0lJgldTFH5HPxXQZD4GB2EdqyinDnR5EM60CvYc/jJp
FjiOSC0R+5+ob06DYDddhGYUQonmTQEa/pLZzEHRqedqWVcJzTk2MjlLGySvgwaq
EIW2jGMMaeG5xv0WvzwoHx01PcQcv7N2ev870ecaeL7xC+ZPIyVlloGls2mlYHNB
bIhRCogrRJKaP1cElBF9n3PfkNCeIMaCq20Ak7NB7LKw2CzJ+a8w/nkv1bIzxEyk
8CLneyUdSs9GDfrMEcohMz11F9TCNs2w8f9LtUhECbG6SXMrIXscYYNvHZjDiJtN
k/GKiwFcQ9vHN3Ro8diPCVypKlOIE4p3mnu7K3BSt0wSwCKuE7rZCVtyFEc4cbdl
uvA8fckopCzKHg3aZQyx/yCIEU7z6TQAILutRP1xRDflqCKa019ZN1xZZyk9m8Nb
dzZ18liETz+FLxZh6d5R3U4z0gpe3Wz1MLwNgNjTzskPW8I7CiMKyeBypwm63hH0
ihtvnUo6FiBjD4QYYljhnqnpGkdPeLf+ajcLlmprZN20H5WIx8khUi6NbxVLJZ03
FWPBmvS60rGXHKTxIq+x6YGkvG+BsVkabW8dDhsxyyDKwv3O8Oiw56sYc7286vvz
2DaKCHQF4J528n/qFtFha1nIH84NdHqhqP/xp8ZD3m60YC3BN0SMeTM48DSlprup
EhvXQKrjuF/a4qxKcOhRDOmYsefrSCcYoJzgCFLeMSRFunqFkI1EyOGGv8ANtyIR
QMdeU7fk+W1Wz0Tm7PnYULYcH5fbDWtK//lU7whWMkrWvGb6XkTKHyPVJ9jgep5q
h7etSsQ/5W1gxrAxOh1xZqcSYPzpcd+kfp+zY0Xwag4i75jZGAs7u+h0hb1YpKmU
X5ftcki5hLs2BgHViV+dJGQC3zZM1r2HVcKf9P3JYZl2HUV1UM2tYgcoX7+JDYLU
3+TJ1O7opHidniIRcX6RggFlsgDcPc0aq2q3GncQKq51mD1VvBdEnZ22R5GM81Aa
gi6VbwjSa2CUPATJ0Iw+UYmBVFQZMTV4cXpn1znZ0De91ubPS1LdR+G9KPMuwOh/
gmgbeQN2yL5p4MDwOwMZryxeFGjVMVVzwWsuGE+VRtzORhqV/LCqbatEyzp2p1cn
KoapzqmCWhGOOXblHDOsAQmtB+O4USLvx7W/eKM8DdLfzh9sfY5SdRrgi/on5nVE
r3hv2qGsNFYbFHehaV6YzwjBNBxbxsa2lq+FydYIRBfvo/93iyf3xKPqhNfNdPvS
I1fOJXGcRqEqcgt84TxH4skOsIayWiSBwK1XKcSv+Zvpp3TsuhClHMrASO7qz2Ce
PxBxsrarW2fZZafyILYca52YY6CRAZw/fOWZU+iRFuw5Rjdtu2+aAZnJZbIIZJEN
ReG+z8B+3hNaa8s0ThksQdJwfKhD/yzekY4/vgu9NmRfEUOtrxyMibR66+OqNNv8
+2HyxpF+i9/YD2GcROA+PasanRmJVqB09yx0sukuj+J/YDT3ktq1MKBgQFKCxR9f
b6vfL5JvMABVCsa5zAfUQcKldEpnGV/pzIcCgt3APvRApbeHp2hIltvY94hbUvIT
ja0Szhu6s7Rqdrwd4FxLuPQfLT+lw2Y1wtIhzWYHw/vcBhKdPsjar+1sjBIxGg4q
yuEEo2eIgyJH5iiaE2CFVRnGK9ldJPrwHOSEXZIN2P02hFzP95f8JSaHdHj6uBvy
neEgytc0VeXj67OgIb27xoieR0X+h5Yfwrn21olKRSRBte2bHwxW3bMrt9cBmlJ2
xVMSxYcbglu2ZHhXyHPRmmMPYNq4PlCC152OAb4hLyzE1ocXBYrFgd+reDxEMjWX
A7yiUScJ6Da7jthH1TyCozVpptze9alQ0B7yI55fQehTmPpzrnMgxyh9KoUJcPTA
N5xZoxIujUkuum/3ihV6gKyXTLOqanMSBBwY/EIB01DU0JOH8KNIeCxkAFvOmfDq
7uFE7sOXlSlaXAeF1iv/rFAhHvrr/6+5mj8ndQjT8QcpINutt9nvNgSfTDfV1bZD
nUZl/Eh8Y//9ipwAHplPcYLFVWMfzJDeNDYsohE/JfptUcawepiNn7vcmeDJOsLa
aKQzRxho6VjlzI6jkw33T8ruat/ekLiQgAK6PGw8gRY60XJ/HpaGIpTN0PwdJY1P
ud1ufXDaFPmEf9ZYTnh8DdUKmiMW/j0uuuG9vvwjedLOsXC5Olt/PlSV2kj6LjkF
/ZblaMEjDIDo/l8n8l4WnPVWuTqBsTSWspmFYRvN69a8x2ScRwONxnqxhIEBiNo+
wZcXBpaD/ZLq50YI5FoQ8ULf9kLm3AZPFlZN/4ONJIj2bfo9LlCnBt2qJGMzW9Hk
47bWMZKOCb86mS8kSwrXtygOLa1ZkPhm+4osx4Ks+dOqrG4smcVlTec2DM8+Ytnk
+3UcSKEVEjrcyVCLa+FP+RKqi7O5BbI30154qefsizskmHlc8z5EVfpbhYiNtmaW
sGtS+8xIxdHc+BuEbpCDR0YZmZNfLdG31AmlR+OjUKrSUMKAYIqcRZ1r6d52YbpH
1XHS5N1AzzUQZGaGgc293qQqSBrNdoLe7/GnVP6tpejAx1mKVcrEJydeaNyclK83
danuYAkYIGwsk6mkFiUkq7410ow9Z6APDMb4WBR4Nov7nkvhfCRodkTPHjF4qDUy
ubA34vweFF/h9UyoO8KKpAOVuI2wqK0PL9FTnnO3tGJDh3bFTaFqsuEdoW/hzWh1
Y3l8jdxDcgxxN6mP+Hn0TBW6gFbZ0CAhd6IHxH73rcJqTgrKw3cONFqyU706/hph
k0Axa5GpWa1vr0eAmF9nJ5VEsf+Y6q9m6iN/FOrJiif4Qisw7mcV6J1hOIhQLLGj
YqFnTRfShIzzsC4jKilsbRYDp5E9UfaZvfldK0k+tuSh7XjMAcdHqhdnR0f78QF9
WN2L7pBPkEbRT066xqKJg8zetexGx7U/JjJXrTlURFZPgNh5PENYqVpLcuF103bH
2xk5ldajL6TR7rPjDgOQB9030pNNnS8td3NDPp66/iZXGWX50V241DePyzkEF4MN
YXjw5TAJS66h7U1yfBF3QGlvU/Hsa9pLrFgJ3Rz4FQeGj83A01NyMj2ztJinq9tj
fZAJ7QNzV7TAgNPd6OhIEkIU5IRbtKeIM5+eBVz9iUTmQkO+pqL09QSTjjnjZLSo
SPOCujAJEj/oe8aIFj4pk0hiYRY4CcpCvbp+YslUiDeURM2+4vBwTPQju7x7PnfU
+Y4C7l4nfxlrlzJAexp35TvtqYZoRpxLrrehnYnYpWYIKJveuXBcMZMS3/lWq2pV
v8HWcrWAh76LohxiyoQ2LZ0bsaoJmiIEOwZHcD8zqr65VfH1p1OO8XCp5RhMCMGe
c67i7DCPybRDnlWIM3oxoBrOu7/6wNWFP+TUvWfD7x+CGX7IdCkze+J/CTyhVnly
2k1sWcYlTpRMqtwZg20nU6rNiikK2Oqb80XydY6R4gv1GcaYHhNObt8BcF95Rz0Q
4EQV46xH89e2l0kcelXFBeitNBknjTyG+WQMP137bjrfVJmH0ZyOd2bb6ya/vFZ/
w02gnB+rJSbQocZihg6PPhkJot+Iqk2HEzyn20QpNwXmkpoSBNgo7q5YwzUy7HA5
TmHRf8a0EtURQ3khef9D78/qAzfNkFZ+t5w3x64kdkD9yomkWe7AWJh4KEae+0PO
ctoBe1bzrBpidE+Xc27RgmQOVAtAWYZ7c5UEmhUHR5uEGYKp7zVpR3NVuRNwJh/Y
NywfRDDl9cSvMuIjXHZT/a1VF8JLk7Mv8DM7RSLhCGh8pJ1fSCx4nE6JYEQG5Dyd
hyyFgYopBEPgXdaMqzQT8vmowwf6TdUpKtddRTYgjB5G8JA0pPDJKmtzPWtgFTG5
ERm1Q2tjGQFLqzCWjzSj8+oyP8UPOrhdPtkul39BQ3MV5s98tkRk8RFhAuDTZZ6C
u/CyxBcY3Dw+NX1LrL2ejrYzNO7QRyFaNlR6GGdZD4fal/7k4X3YUTODwpMzb0Ag
Z4VO4fvQWrisfRqcYRAcHilSfUYGARODAM49Beznw3ALSXtncZMMdbOSXIOQLVxU
4UVGpO5It70o7MNobc6nIfzMXOOnfd2GEU3pdVYI5vtjy4kyv2TNWZHhgPijH6kK
pXPWePgC+ujlVJA+icl9bhWYMFQPSMlbTm8kiInxoRlchIA4cgr5Zq+gtP4XV03P
YPlAm+u5JXFLDeQIk7vH30voA3p6NW1vKjgKMTOMX4mQY0zE0wwcOtAE7xG7mnoB
3Z6dbdGQTGgeYia/+3pYqNeUR6tbBYIng/Laq8Iq5Ft9d8/dTYC2FJbpp9tdJw7Z
F4/YPpYHYUE7FYNgCVXryh+FIdSN+JIhVkDO2up+vr90z4B2GCEWWNtz511LGJMZ
czuqYaAj0Cnaw3n5V6yMz6ChfYT3CmmeaK1+wUTi0x82v/gmrrjdETb9wZnoMYV9
RLBeCW6TNvdr+jUdOJ6H5g3FtkeBvrQs/Y7NBU30xyTJT9df04ofv1c8AY+Dyn7z
tU1N945L0p7WUmavgW2V2Ul1yNesEpwRpQ0no0ZtSDHM0K01l8icK9twSN/YyHL6
tdlSIKQsB5ljYdsWQGCdbgPHekYMFzwgURHgDpSEOkytg88W6p1He4nAQkNRt/kw
6yIb+7KcQ5tOOL4eosNaF3s1MPlzF0Pgja6mduGZcz7dGc/hKYWF5SfvA3FNa4cb
NRtMQTY+BZBw2krziFfkgvmBbUOQ6YCEDHR6DYQjCVXxiCK1GakGlmkMNZwUTZev
DFaHHsxIvuFBMgl6kPKB18sn00kr7j5ba0MSLef4kIWJkKiMuQn4dR4nzdOHF/V5
wL6RVDlErfd/ZbiVElHzIB/5UtgIwE2i0xxFbIfhpIOlkDMWnNwm8hDNUbLtdl64
75Zhy2rvLB/lMWY5Xv/EF7Nu179tgDPXebmULNfnMRPce147w2Mq34165iKvPto7
N+5X3vqAjnyb230C4K/egms2yN0pvMhdtDIxBUcpXYHGbPwBpE4Mu+uWD1Sc4MA5
djwW2mIGRGya12IozSmBDNSJzpF6MpLOdP/ed1uqcVNvETet1W0B0tyd12bCdYBt
/gla+7CqFmC007ewkwgFSS0FrlJD31XJ+2yGyeYgcGedMlY8rurhVaVCnlTwblsl
UME34/khC1QFz0N1opzHIhuyr1AVWZmrTxBMGufg20Q22Jd5kKfeNntj46GvVZbh
VlLSf8OW8alaxp7fRDqLWbrwfE+hrBwfxJ866E0n62BjmlwIgO6MHarb3iVXn876
58CmopSmt/oCdKyQ2kcFlrhBLnDeeCfWDH2Ovw+SpN8thNWuniXe4xUrjTx1gFqy
4NV2PHSAwArjvv86T2tjREyUf5Q8kM8McaEnMXvLVbzv01VsEBcI1mEvlxQk/314
+Xj6xlJDynIFY1eSZC4c35ILsF0I78ET2Ps5Ks4uhAvKevWLZsF8mf0Q/I/lCs9x
3eShpbmk/yq48l83A8ERL7ypgrneyBUQOXD65IvnF4bjPdOKcmrOI/Wbdua9OV1V
HqPbn/iwjV47Y8RlMhvCs9v8ye1o9gt/t+cW20Tq7BiLkhNVOafYzYnZT3ZAjnII
ogd30oA0dEEeajINY+z1lN6ccBT/B+4NJfG83jb+/B/fp3IzMV/TV1G3ugpwAkhT
QhrXHAompAD8zHz/39hKxXwp1QoOMxtclb3KqVkDfOPobfm6UY6At8Y30M11MA3z
33ihNMRuFs2PAVZjwxjwuIxvouJ8Z/bSB7mW/TJZ4Gt3LD2C/uaBLeDRmGBVpzgR
EwhTFXCe5v9dGiyCW/8aNQL9FIgRllJZRNErIotjrOqYIpsA/Yfah3yD0iu3yG8E
2QP/Fz0CFLWr298v1OhRpVI72UK4vJdt6QZ1URwvpHbAdedHeLuN1UNdPYiH4MbT
M3Z1U8YnIm/oAicmsNUgVLvId4kGEE8YQLdCNize5HQHo1/DVSjOoylpqzakp3w0
6/6CoNCmQiE9e6wi/CQ/NOdRjPpLlRahamuFFVB8lhuvmHfh2X//oPRhsInaklO3
cmujOcBhoyi9v10b+5qCihj/YXiZhExK63QSO1aD0Y3j/aiO1QRK8MbznwxTV/Fl
7msjjNyAkEPB0HoGrZvwWtADxkKAmIGIuQiaLJTSwNjld6+wCMY9lCfA64pNyFsL
N1Opjma8N4JlgUibriqAINi2wVV03Hoa0+bBQEVUstEyL5UrVAOINM3iRh1oebWy
DwPF+FYW2XEa7UA5DDjge2lCcDKdfuAubGjZ7f7R8NG2UKamzy7XTm2KLrmcuEo/
1wu1hMlJcBN4UEDD/S9yV86qvIfD9otMqbg79+8BLeQriFC/7t1alNOgmKPWMWXN
9I5W8ZzFq0AjkDfGR8T/s1VtIhPftC0GOZL6XizXQT1UhatTP6aAf0LcNUKvIYfA
nywmFlCmhFV8pizl5usa6/OJG/XjglyBMlCmZITFkNQV+iE7t17WI+mJu2c6kKOA
7/LQj61uq0+LBzoDQ/LMOQvGN3A6SICs/WRFtRHdRpyNoipW5djUlwbiSVjwbwXN
EbroshkBdMuRZOkxvDkMDbNC4Sta+1d1q2uB0U3G0HLB3s7t3D/K2zTLXtwHprN7
brR+2mOkq2q9oDn/zYCe1//nCudSp+vhbeS6Cwrch4Trr44IJ20sWbSbcfdnzDnE
vE/9YOTZSCCSH8Li7SwJ/loghx5OpVP89doD59o+mGXRh+Jyv/SDUiWyvjFIh0/5
tiHDmM6oCFktgNghT7Q/+BZpDwCJq8cpXbavL502O14SWEK2tgEdHY9cCgmG6jVe
SzmiK2T4waxlykGpCqnjtDI/U7e+Hky+tG8wAgvEGLCP6olsH7gLUXQ1E6lARSuS
K5mXpWNmYjGtb6jiBOCHvmuzZF1xgmIOYZE+LyLFbxGILOLWfW4aoxgEUNdNZsya
U/SKdop7mkF7PEEG4A4zCZVzW2TzBclPz0EgSWqNBI+eAH3zDfZ6tWCm4ePVw57P
aIAM5QXOPrsWmBQTsXd1hQFD6nQVF91JaGhKS+kB+hiYMtbFwwipEaBACcaZKHie
Qp5/EQcGZ652BXtVp38EjswFpAXFP4PUjn9ZC/cUBr6UotYXnH4LGtsdvRV4/XrA
sIYGWNafQMSwLBOnUQJNjy3BWHBUX/LP5WcLsZbPVKHm1t3CeS2LnBxA4Ir5ZXVp
Z96EllCXnaMQDE40dMz5gmUoSOpH5anhPmR3AYLrxxbODhIcY6kzU2stqNVmVBKS
uou4Tgb9Nh2ZkgIPSUO5ErhCF3U+A1eNRkJVHz2xcarrTCWPZAOYse7YNu2nKERn
zVGIOWEzmL7CFvxi6e5STUMUdMqKh5ZhrL1it8GZppD4PWdHWH2RM6Kdv2yTWFg9
k5lk0bVwwEwSq4FnDXmcBVAXBRymK6QPCgrrSZBCrX0x/TjrxhhIQ6Ok7dLVGvj/
t4ir9FWGBP9YnBzFC2Cx0pHui9N0HJyxfKmDZYDIFPwJR5qrBIaR+DB6i9L2r8HX
C//CvoAzjIl/ICiHw12ghfCKoUSZJJiKZJxR1WPN9WZ3I/SJKcUZMKx/VRZjnreP
0CGnnwm81MohzDK03fBPsn6lOh/3041xFmG4y0a4YuCLlO7L0ogVjTPX5V9V6Bv7
pqeK4oFKUUUoRgTVKgJaTzd78u41nl+Fj5bH7s1pPAT6RyvbF+RpRzcswf52bfhv
DXyEX0d27+GjODfYcleVVG78GA0z40twKtPzWaCz7HIFzQF3V6OLgt7DvrZa71Gy
eQ4DndT1tg7T5+XdcMHVyvhto6k7bOLLt85H00If3SwtH7qtHiooAHIDymtvjzXB
+6VpbNRgR03H7wnk7Ik0tgh5Qjbmf2MhDBG4z1fJOqJzgNH4kdbv33dQHaOxfIHD
zsQSkh254gTr8Zgt6GHkEXepIpG9tE5iU5bQRsPmnzRi0c+I/ZEye5gu5VWDQjaE
k+vbYE25eBcbFNmsecR8UWyIP/kNdzjCSZZtydOqfmkM46utG2S6JGo+AJdOVcf7
Tzo4U8ARsZJ75406JVCWZaTO9+Bl29Kc2f+a/7F1dHfV0tDRylnIW2RgoP7CjVpi
fZgmzl7Tt7XOawsO3VzhaRvMZFnOSsy/f9ieNcAcZFpaZrAuDyjlHAHXTGCLyzMb
ASOwPe9ZsB6PfksnvUZyIdZSPCAjBjXQv5gS2oHT9VNM5qWC3RSDSOy/t2O1uqZW
s26rNH5K1ji74lzl1fAWkUQqkl5DcM1RKOwm5iOnuqFT9PSs6m3cnXVCTvjNFxyd
a/+NlmdoqOBBBKfSUEFgLN404U5F2SiggYznQbdS/KobhkJe6RXbWyaFGJBdUneQ
xoWkP/DkZt/aqECdPTWuADrdWp8MQH4wsQSUwpHpPB5jVuO5kQab+PqE9PW3cewS
2qymwno2GKVBFoaSSUJPn8OWkw4mLCo5zpHkKA/1Q2of+m8cQEQHWVV8jzNhbzKn
qvf2q7PjoI3fdzHTNR1UJDNEhr2pZRN/3uJmIaYwgWY6lAAdQS3BRY0Yj42ZTuXh
S66kCt945OfHq7YL/q7vhZdXw7vaPS/hPXKbSA1ye163FQW9M5x0XVER8v7aJwfI
irZH+GZ3LZa5a3SOJWxFnvwuKHtNPAu5FU9NE2F/IrvKKUFAsfKaiBTcn5NIKKtJ
m0oVHfQZuWxM/1F8ug+50vV28JwimhLQepbLM3A2o8G660wWF6jHAe1jS0RdQ2PO
ylk2ezEOzRfseRDuNvC3oxiOfHP7+v4mFJ+nz5eltylVCouL83dnC8aj/X6tYRYW
zk+CzDLSpClXp2lfvuNBz0dZPHaz5qpoMbxdpEhjZ1ZLXeHSo1HwoiCTYj73S+Mk
Zp1/c/mxTqXr3fv8tLZIR1eGPoFIexo3i28nrx4aRIWHFJ6z7JLVzG9Ecxmd/dUB
GtxOaYuBj/LCeAbZ6S3ofd5R4oxNlwRsjj3rzSK9KVfDsCIbyU1PmEfm8bBGA2kk
OEqhSLLZztKXbUCdkuni+iypXnntIpl3qVF03dhdqdHW9p7dmGC4j0YnXp/jkllI
g6K0cppBWFkyxrLbrPqPgGynnkGmauFRxKYGo3WU1ha0N8PwiPfO2ORd2+F81Cuo
O0TODV7R8i4LqsE9KyD4yQ3OYkKhKVAeiIdRm5imBxe8uYVIqsH/qknnyGuwzKVa
OdXisNN/zhVZpa5ek0Fr2Bg4vOrjcxKTIeJHQSRrv65F+bukonGo/drVKOjdJI6x
bN7M7oxEdRLqJmwiDm05zBUxt2yRerpMBsZHQG/rMa6/o9ubYVi80AIPKzDyEdAa
qwvnSSj01ErgRFFpeeRDIIrxS/1y2cX6feQrNfJk2CLocaurV+kJD4EmGnAVl/ai
7Syma56LLfsRKMkl2+OBuAhnfQHZ9LfirrfUyNdzhrz6mUiAty+2KOQ8tX2PFgs9
DEYQI9wn1k5x/p4h+lY0yqBYgcaVKzZPBo3zeDn3OkPEWMfNK/BOcmJmp7Pgg72m
tSPWLU1wuIRWXO3PiDexeViFsaVtfqj/zyGZ/Enwe9Kd1j5Lu3zU31lPjkmfFrf/
0P5ujvaswVMCMombv9g2a3jfua5N+z0ECUGAfTxBzWwv1f8DSCLtzpHYhsBjH8eq
1us8kxF6sAOOyN8c0wBKPCV3PAXPtm3PUcvoETl3m9SEzaHfZFMoCo6eeftu05oi
AeXPPNBeQU2OcH/T0AZkI+unygXz2c84R87SCre1XaItBlfgGZdC4sbFs46XFdRz
nZk7zOjw6kEopg/X5LHu9FG8qAccxwWem/DL4V6Jbt1ScBArqt0RgwC/+h4XtkSn
7Q6HsGz+YXgRMqg+5f5Zcf1WhmOHBP4zcL6ohmRWXU+QzYKAg591E4Z91afmt01y
TkaX3aYi+UxZDweVA+fj3VhQ9DdoE9+UYJpKdHv6OBxaX0NFGs0yEeQnWV++/SaI
XlLyXAkqf2zX2HbOJsCmQn1zdiLdeTeb0sedYHW9bN0xVtoBO90zCw6t/usKNpHA
Rizn/D6WrbFFa34+x30gJNtSsX0mPv4iTY6UhzgvEsW76Uj9ABe97urPC35debwj
zCeuyEnXeAah5pMIjq4w5z/dWPAY5mE9QVmfHNVU/s6A4PfeVLBV7+HRappAeG+N
BIYghLe97Kj1CklF87p2OnHPsS4ySBPUZNqIduW8vRgvcNznj9CHwdGDEr0WTnJl
bzIUy4ZINIS2wIjvZY55PAuPxrM4Abw7x97BEspOYCuQeq72b1nk6GsOVM1LMGu+
TR0lRbAoQw5fJjMt/sH9P/aTkf6N2ltUf998ZB1AgzbiyBfCKcuPKG3KcSPpUTML
AJ3YPx/G3DLFjxo+M8W0IY4rtWePMHZKPqYluHv951Q9TRDggtNQtQT6LDjdDZug
A9/2mSCI7oAfml36+93gu+G2wONWzWVXAveT5BOK36s7Ooc7qVzV7Pc8g7SAMq1p
x7+L8Hcslo83toxY0WMw2Eyv7d7YCzWT+pJ99ugAU3vJBytRmcjZrithUb0PvRJY
ogVzMKmPC8IaOiJLBeD+KzvP13NkW8vkieNQLcGhFw5E3LuYKDG11V0J6PfIqH6O
RvOfwT1PzBhY4OYktPh1vVzZNauLqAWwYhKa+LYBzjKMalvP4sw3sBnL/xkYsL2y
FC/K4KaQPx/ftgeucITRVzVSxUY/cYcQm5pLQlRWxoa1OC1c/q/v95ETBtBJ5qVr
sJK+0XcEtpFqiDIz6bbXB2OFyGZimHDE4aH5DLvY/XnhJI6aPMLOL3EreQlz1b8G
Gxo+5gFy3k6x71k1pP5CO8JC25i2cRM976rSX3EMS3WcFZKPYUDd3cNxPDzVir2I
UK7Sl2VRAgW5tpEv/1DzodExJVMwA7HcxP1csY+Lp6EwnwmlQL4wEqsrLkn+wtyC
70AdMsob6mr2GTmtYlL99oNd2y1qke5LoheIqk1zi0DzJ8lSB/Wjd2HtupY5k+6o
YzU809HPRJZeSB+O1vcVQyTysMXuECMsuhw6AtYCHn7RD4adGgFaRvu4yEaQlnz5
UZ326TTcRGlfhVeIKFNgvjMY1KzKdHM8HKmU+8XUflBAnNgPq79K+MFUv5inZiE8
UMpe8PQMwxu0FAEMHwjwU2RNFXIRNkZlyjhrz3ayiHFC4bBAcNnxyL5zxFxm8hhJ
+ONMSMHkum79vJBXKgeytFshWIvv08eqQbITx11p7OIL9bDFdaWu0k+pA0oJ7r/o
0hSqAP5Lkaapu+zmP0bRFTAmlu9drT2ZlxTdTD4Yr9/EDaXnHNGW8XS+c4qWOEVS
b+d6UhUHXb6rnho3UOvdZtkUnnvJ+ptzfUUw1RLb/4OWZjaAzYnDVwmH17OmHViK
gkTqK7PR8c9o5EOT4v6Koq/WBGzE1pLPwEdJ9bYPEtQpX36Fes2m4sIt3pJqtyIp
rzOD+lgP6QRhHMObLW+FRTF8axmA00ShRqNMIlqOmaN0prWjL1/Y3o40yske4QOg
1D+EVZ9Ee3HyjdTUv9o3pSpmwRNAnKVMy2kZK8MxhaZ+5heb2hjwe1fTRNCPQ2TZ
11GjhSBcuml4zKNwmPCJKN764s3DK6Zf53zZA5cs0SGfr33TiQ+xrxgnimJjypOP
Y+MdFwY0cuDtGifZfk8kCSqVeW6i3++8AMLpYVk47cwbQP1m2pCaZjr6H/3iUy5s
ZENxsUSs00cqxANvzUZ1gjuehjSjfkRvI+xaa1b/YAxDs1xBZrctIUuOLvxnZV1I
Qbl80FYVRVLed0Ur8yhGQoOkLI7pS8MWa7A/EwO/mQ/5sZ0X5SrQ7GG4n2RmmZyJ
28fkuQB3fN6dDiAQy6L4jLdtsSSgN+MAfbMuKs7GMm8m5kSP5+y45+KOD+gVnQYR
GvSTxyHT0kVz+PEh5XZYn7vnBcXCPgVwVJjIxOHFn6z1oRscGYUbxD+r2BRov2pk
+lxcgd1iXQU0M34KoSs8yA+hTxT7lW8oY1+lpHbzOwIv8/VY+dhe/K4ZUCDWyPxG
foryK1QX7Dp9QTXMiQm/41IpbQPmgLxybfWgcWjs8FryPtPAnZVHIcWUey9Hl8Ni
L9Ok8t8oJVpI3GUQFfx9+PtBn2O/XqNbH+qv+ov6FW9rG/JpF3YARG0XeGg1ISCL
R562YBFkf3GkUAVjTfbWJpXEvkN4c11/HVLQxSBvyJ9GBwtYNZeJk0jnW6IGbU03
BzU5L5LFleqBSEDpSEi2ANoIX620NLa0PxNJ2oGH3HbT0yufCTM0yu2i30Fd8LVv
D4ZlLQVSsI/3IEB3q7jihT5IlsWIenL0bbDFTc1kr+xVwIp1C9dIdTjaQE47gNft
vxu5DJLf0gD/kHwNLyA7qZ+OiUXlqBNYdeYVpeHzTF608RgY8QL1n+wbQc8kXk+p
xXx2B9aPn2ggsjD8f7ipLfkG6klxY1VZA+MrUCgLocpIsHfDjLDxpgILUy3a3MAi
fKuXHT+PLYgWara9jdcqB2BT8f+xg4Sn8y+EOoy2cvnVuKHeT7wcurzmNtHuub21
y8n9g07/8eGSiJrbAgqwsF+JyG72AD8KINq/3rGH9TJibuLTTpfSmAZa6k+A9KsG
fwm01Lyj8zD49NIMiiEBbR+txgm9n2tf6UiVGc1EzRER5Rk0xEXQ1SfnZl7091Ty
j/nOejNVSjZmjWg2f25NqCisI2oMxgEo957wvktZSj9sx8xqnhJU7nnuRnuhXfJ5
ABOp3gnj8fp7NMb+333h6iwoI+yi3KoJQYWIKpG3icc6fAG8pWJl2W7HQ63o5JV/
sIHFq1lSjk4+DEXD8iXj45zkGoqDklTBkSctvt5PUPfK/BKnRy3zaZUnmDD3kzuA
/yX5PjNhFMM29g1XocDe4edEleGkv7yLH/WTgTJf3oqJsSN/PqPgaWsFtu6vx0n9
sahr3FlEDyVHn6pOs310XS1z44MudVWqb2t5kuss6GkMdJMmAt1DEEeOhvvEqWM2
C0Q+BzO3Z/qxddZ2rksSS3pLyLOwzOb3PC4u1chjOJlRAuIN8pyHmp+VjsbLIGui
Nrfw9o7fMFllbJZe/+FuudikjT3WX1F2dum/CaeOmcAJdWZnG9etWKsH3hyYEVbY
jmAeFkP6w35VLEiTf/H+UFrSZQTBXYY9aZ1uLIhhBMWTzoF0fiyGB4Du42XnudqB
C0Xj7IStT9HWe1tNlCgNCbkU7RQbaHIWWJ9aQpVXpC2GByh6UzlmCCthjwEyeOyr
kSgRUQVvIU2SIEw/tZT7HcKPX3kMR4u5FovDSA3uMeioMUZv8rOXQZXW8MUnl2na
RcGp81+Hh6k6kBYT64SxYP7fGKqtwEDHsD4Dt1fTV7QJJrXK8Zs1k34HSxM/X9dz
MmeEhp43zxJXEwAdApwvl6J7zXM3XgZm/DChSeyUwCIDgfLIiP8rW4av3D6C5VQN
xJDFy7M+0FN/+Nz/QG7i2fqJDeAQXcOiCudslF1JRgEOLsr2EJj22QuMnltu3rMY
sHISOql8Fd0l4AW3n/dqCye/GaVLSlGS8u8JHOO7lz80e/ThYw9kaU6zh5+QuXAd
aIGfxGcWZyR5aKLhBvuS0yfmS686DEKJp4Fb4/q09Up1oX3MmBX5OZ4si3UwOEIp
Xz0xnvnqi+ddBG4Jurb8B/fMep2QOgmZ43TirTfqEG8s+XHx3TARi56ZTyK+ct6z
3p68vkhJ7q36C88zEl8zqvpZo8IRn/OpXV9bt72wAbzbo0Up5eyaZ4gJb7gil29M
SJac+JxeX1FmeiDKxyer06nrEP331BNNm3HWzdQuHDkt3tkdq0dAG/Re+2DBFJlG
xmeBv6UvLe81JuUm8Apb+CfjuQTMy0OWp/G0SCWDEeK45hDqUszZSdFPnLKqDbCC
84MDiH0m979tLcKhM1Zj35cgtg4lB8E18C14qWIqChyrTALuCym02GB5pVXvpoBg
XLmMQOd0Tansg09RJZgl20ytVprqQxwzyLIb1iIFJIn/abn1vfWS9GrlhIT6GHW3
a0kdp/LMWraUP9NJZiZcP2U7Djv2U9CEPALY1UCR9NZ9FkSHUAG70qjhiMXn6Pq6
m/uvRQq6FDbx2ZdgXO+qTQ/ZYPUVclOvT04nxnjGC+xTBWf0YKXtnRbFSokl6Khl
YHj8WLZWxbVHuoDxFs4qavLTMUrWlj9sdaWYUXVBLBeOw1OlviMGEc9kjTrurP7z
XcXpaFNMIscdYMkewZVw9UsJoZDrxpNo4z7i8d8EsAdckxjvvSgAAKmgEOEQr8Uj
lr4CTcj9myyxideE/ZyLbxScwfIaDvXR/9lrzRD6MNq54XGUzYo1X0yQXZE9apJz
/gnicmStd/JmMj9ffgZo84W0irkM0cyagjfhL50mCySTZuiQXMh9WofXhigRS9cI
ZjQSAmy86tEKqIucuu8ROdAbq570PmfodVGQp55jVSsnCh1gBq3DrAhRidRXio56
H2LlWAK0jpCS/pVd2Do33i3O9TvLNhEXpVbMzZUg46LhNUyph4ARqhq9oNQ+Nxxd
HOVY8e6HotaUVMNR1MG7MVEk209liyCuFzofdO8u7O9NCWZodvc75vHixNHSQwoU
T/dvAczwVR1Yi/8kbETPOA8Dl1UDmgTj95GNU0WHDGrpMub06CA8Q16yY7Z0+wiq
afnVXGbGXrjpC0bJML55bRweXk7OH80aPcoXZ8WJJOx3FC+jOi9DKY4i1HozM0x2
YtwnXBD7+m6aEaAek7QfkaAMnQCNlhKSaDPMCGLNIFXL7l9oOu2UMOJlaqqWm1XA
1JJQJGqpN5T0qy7QHHHpi2IdRMixGPGy6A4bNXLSzgUs1/eSO/EJOGBN941+1Y63
OFs4F78aaxk3FP5mxwaZjOFNghPyr1JreL0V3Zgt6+0fMfvoeMnpBhu+mVfOXf1R
X2GcTM+yuwmYg5T/xXnbhefp00anDcLJZ6SxSLghvfYpqI8HMoMjhiT3705d4yT+
LLcs2segYAjLU2VNCESmJcS0PhvqTPUhwnnRrthzZbcW5u70cle9zZjCg2DlyaEa
Px9Ba30JOlAg3mza6Hn3NdPcN4uRXB/jRbQp8F4AWM4rvekNb6TBMN/AOQtgR0QP
vRrHQfDurDhwrd6nZ+ViJrN7iiQsnAZpnwVaeX53wiu7aoGpA63T/kD8AuBudFcv
FuQbqmoZQyl5NEpjaaxbjPN/nDlMX4FSA9E/sz3TAg5JmDHFkcLb2VKY6iu5K9MZ
qUsmbnV83R9tC4q+tRpUskwUWtq4oCG0orPVGWtUsCb2HBc7ploImrZOjt6fFQ8i
H8w57JwLuQF5wREhZFphZrE9+B1HClJSCK/jBDeHIDngalkM0SlpgAyKzuyCdfbl
3GFzT/N6uK+bPgp0JEr8Bp4gcfllvom1BVuavtMqu+UaTJkPLnS0bp4eRSkH2Ju7
pigZ2DKLNJJg3jBE9IaAOqEKydjMqoG+Fz/cTN/+b5SiLBS6lNQxENK1bv4RTt9X
49KQR5hEhGw3O+l08ceC3oVvdeQ1ZryCMwvNWdZ8yM6vwm7PtVhAhWPBAo32C0nO
FDByy2UcBQI8VLnDHurpo49w04FTrPk9003VOFyFvo2GhAWftHzaY2FEY86y5U6V
YDki4JzEbFZXwSwVYw3afSITOH0wJzddfEU9S7RveHb/gYCxgR+c4AuZ/hzeiM3c
0dJ/HElpSVDifKkgjS+XlVR3bZeeaAvJVfivBUXqNHamkVS3s5fjb3Tm418l1LWV
Z7XbUaVpmucEogvoYDisSmP87jT5FP+HeZe4JwE+ZF/xr1tkO8f/W3eARiOJM9fr
9gxFfve1FUpG9bNMSmtWv7dUk+Jxzy7nx4NwR9uOHoY8FoM2/0sUPt/t9P6gl6kv
30mVWUbC/9aWYFjvQWT7ZyMftQny3crS/H8Up77f3VjOqJWBuCbkc8ROdzaYmuK5
BEXbGXgh2bI/GNOkYAOzeRRKGpDtvBmis3vBfsdFb5P5XXMCGSDV/HhwwnNqWURO
uuSgOT6BNeXpLuK0GdbjUJU5F8NoOFIDOB06irgDhjZDDQKF1R+0vfu1CW/XIR7M
XhdDssx9tHk93wJlKyOUOJJcCP3MPTKDqh7nTrrR8gKSjsqj+3a4QQtskKZXSgVJ
nMc8cW/I305G+myansPE4wVnuv2OGj5qfWZdEyu0BzBo5O+k3/pT7oIckte6K53A
fYWFHh416qcIF0C9d/ht0riFcAw/GKje3wBJpAhellNeI//fE8/eIACEzPOxwd3R
1S7+8VZ+TeUUEWnjn71ixXkKfgC5TCmvfnh60jGE1jO+Z4OPAVLTWDP7DlfBbeEm
Tuyzmd+uqZ+yCyyJMbdufjF4zK5PZ3qKxsCJX41yclnu+112pdpgrQh6U4vt8/ij
Y0D6YcHbG+skmYv400ZW8MjPHugh3jPw9F7CDJXvx30SYoPsbCAwfRIXGl+I5Jmb
jIBjbQFwJMyux49oVtC2GvMloNGHbaANPTHQoUB5cKZACfATf06zvxxbynlsTdwd
3XjRvrE2LNKwCzjOHkLHBBdBy/VGBCgyYln+SQUAQAwNdN6fjNDT+RHFBNRnTkkD
qhDE1iwzWaMHsHEsLHhsz6ZfWTL2fyrmstNyXe+XCQOPTgeNTaSlcWtKfYMfemt5
XMJ2gdGBpA60qQOqGmQ1adJcYb5qeEvuBQr7RLEajdsiDuRfge+15r75pPxiDABX
0vOuzItsOFPMZC98eRzQWTS5mfTiBAD5pzG4GAEPkkDFyXs3ShxVGn4oczk8o23H
MWituArecQ+MxDGi9PSAfpcQIIjwh7yckH9zMTAs3R6wkaAAcfcdqLfrSLX232oU
j5mUByteI5zhmu23R4LvVjuJh8r7rtxOZkscwJ2wDLXl0kqv49TYvpirm0zZEAWF
851QUPw8s2jKcqEyem5AIJ5medyXldklFjHjPphzRObpThZ7T675m2v+HKkjgEwc
dfqtJRMSlSRFCOjstPk2qw8wn6A/xunXNciRVJaP8XFHVlX7hOX0g9synvIYmu68
dzWzo9QCVEZy/X/YfgUnR0j6hYPjnUqUYSMoA/Of/WLLFbUvMGaS0hs/82YIraTe
kq0y+J21E4dtLvzb00b6CNl9G0sTtqmfmWa//HXefK+5oaUJkpGfOq9aTjYSbfwn
2lxv9XqTPbCUHJBG+FqR/pLJsq9GObsODDXl9znFwzE+UukHGqf5w+Tt3B0lbgX5
+N3/jk4rRCeS1mnHBI87i/VkPbxMB2gsoWkClBcTWeDsVYOvsEwRJhxYXGQaYodB
yvnLClR/IeJGyyBV8XRlPssl6LVDYSOBceV7gR/uQMVSANYqcy0sFiyzJAaUe1W5
Xyso6LqAs5aRpW3kbIuA+Rsd0C+C2S2Myigsjt8DTjmGhlEOvGBhG1GQZULdC2WF
Q9WgMHE248J919QT6MSX0z6aSDX2huiP100E1L0CACeBp/UyGNV40VgzuflQkiSO
SRZeI1ci2XscUbFIXIh0wwBIFtLYSU+AEPK4wxySHdERqn7QSgzUT5BGaOoQ/2oU
3MJ8e0wbd9psg2RAAvE/qvF8EyIevuRd4gnZJUVL6li7OsHIyq5+yOQGx6nvb7ei
csgb7qqXhHBvn/oYi3D4C8yFzD2k5pSw0fjcBC2w5s49+a3P1z9e0Wg77s9ctIPc
OLHD7u1vhjh7CLeTmghlNgGjofsd7QtGbesNEplgqc3+dC0r/SbU2J4ixXLXKpit
WFzhnvNOzvbRHAbol+58hHApkiEOU+Y0zA4xgw9xARAOmBGiC4qusPe2gfXWx8pK
HyrwTdBiroQDzMyqwX4usY9h8dNZrFRUeW9G7ft/COjbO30CmMxTMuno5rOe1+3b
AMaedM+zZDU0B5+U9ClJLieh8oBkA6CPV+WywrQz+UVo2au/zaGm73PxFaazdxDs
PWG5AkbkFahfDK9fBvjZhw/pAq9/9bieHpmZsbUCruvbt/0xXg+WTApFESQu2yr6
mXGNiNJyqTuQjO8hgKg+thZTEZys6Dn+1cxs6tgMkTVyp9oLg8wbf2cSir7p1AFm
fbay0DAKNc/5eIIWzH1iNA3Ybag57O5vl3d6pFk/cAe+OXt3G6C9pU/iNzQBUgJb
Cucvw440etcUZXo6U31LRX7ZM6uNCTmsOZJATIFdoZUIC4AVIYO0qP6jEz2sKOVU
zoUfpFL/KfwZCSF3fosZWx10616BmbaHm4/5AvT6rCRbCbThYbY5cIEdtGFbRQZS
2CxXnO/S78aI5zT7lVBcA8R89l9Vy6SJ7hZ826Sh59UFT2kmCKqKWX3k8NlY33o3
Cyio48/IWEcOHRJbidO6BUA+xjJ8MSPwgjmK2kBykfNelEkodql/+cUPxGX/GXZ+
pH6ajCCE5MZxZc4k21Mhp7ORX3DiytoQyOKqA0t/zKpEwy8Jpg9d6STLLNQkaF6G
r4ch2FevABI2T94AJwjcnse2jEG+d3XsVByI8ls5PQSXIJ5Hhd0Eofz8+1FDaRK0
rJZAyZjons4YIqOmBSHAJS98l5p0R3SF5WEnjt8Ivp8YdWV5ygktXOTKOHqk8CZ1
ahjXenneQA4I9bI7BS3TtNm3NRIJPWZa663JgN5j4g+LsPg/VysiUzjD7bHSv4p/
Ko5YXSQYmM3dWBex7ewaXd8WWeM4+WUYXjl/VAGO+vxWzVjf0hvdCYh4OR8BLVk+
psjdzeOvyGJK2dpyd2q+zGjfGX9NEWgsUOCSgEYYwquTKAeeEcDppcFY0LoaRwVz
6UKV20M3Jk69/FaB0D8rPKshR8nS+IhGInZNwJIvekDmTwosP3JmSh1/wSR4FPRO
WJkEEz2OgPvTIZ1owM0upKxxKG2VmpjgJqlOm9qtIP0gWt4tAAQqlInogj7w+cNr
bu1SikiUKhqxxssR+UtcYdBa7tsoByoIEaLVofxNgARfXs2cOgMxFgR+rcERYPjV
Iq5cyMUwKJ1CeJvICPV16dODg76Ba7RIGd0tmpoksAlemd4novRtQteHaxC5HrHk
B3MatV9WFr1vPqxjxTtMPcG6IS2rNNHLxyZlzrBTicreddNW0nk+Yt6XIdu8popO
xkjzC71g6nqIYgIUh1BvWjfbHz60x8QdUd3KhZBX1bsB7Go3H1QAcUI/13mPcvOG
SA7YacG2gwg8dZzZKZlzjizZJm2QpGUYeHmOR+RSJ/06bjAi2/7PK1RfLK8z500g
9LPFB3HIej8zAaHXh/HJ7I94SopudkEj2JFtlLpq0qqyCOcLFKtThGaj8qj54hdb
2OqQjv51onPi5DllF0wYyUXZOy/d1J/8tlLQH9w4YPc45YD3tdh+YMoZJAn02/Vi
QsHPyBv9FupJmO3USCpXeeBsIxSeGwyPp7eINAUu6Va01wNfUNoZ1H9Bm/QtpRPO
EzLYvHCVGs1MIGNSNeKl+/9G8FjXZalYZm1bLCfypl0HlYqjbyldsZxNwmswbjOA
YJ53aTXdyC6uh870RPzqPy/szPxO4VGPFaKmP1+DYtqkJNnOnFU+6/ASsxkES2rq
+XrlcfTIG31S7PcureaaTDhT/1lC/5EGnvqzHfknM2+L8k9hgNPeTVri5QRn1+em
PDnMgPJCkZkDA8Ahoc4GRSef/odY22YwScuFjJ9fuQ1I2GNkBqGV7S82dVSlRxqf
9OIL7ZTbA3FD4L4ZgCxo+gtqkj9D+h2bnnAkV5JktsTS+1c6UqSa4us8zAVSa2FC
FltOuPcfv/TuHg+59MUeJKb945Oovni2LrjgujPJD87ao5LwfUtgNGOkxn56Wkgt
sezzsiXjObx9oTpXz69XPuRLU5NobBfME5LWao5LIroGBznIjcWqyVd7lL4Ig9oJ
QFmodmV3+f9rpzKmycrPfXepfFlf1+SNuW5xs6tK7ZeBI48xfsT4Q+Ui/S2sXABg
ObVkDEABmYiWq6IxQY5lHS9f5tza0DjHP7joc4D1JMPzY4CQo0CItpqPvobNbHap
qN0LAbDajj9WsmDj8VImuURKFSU5awXzXAXDejzTzXYPmVBG3DS5YZDS1FUCiBbV
SkypZr1VJm9KUIeeGs+dSnRoELWoVfljW0OifYYvrIwrsowzvAlkds33iTlsgPqo
J8HzYLnv0s40U45IWI/tGyG8aITsOQB4ZCJeHWIT8k3DlSaxYuumDAlSPgFejbFo
MFrlbI9aAGzG4JWmAicOoKCsMfav6/95ch+Aeq4NQLWtmUgenCY09XfSKLS/dZ9O
5NsOC+hUw+yapmsj9nVLg/I8MQDExM9tNEr7LE4sKmLUfSbI5/fz8Ah8SroxwIST
mTAGBMhzhrBIegeILJRJG0AVY17ntomWKJBvSvKiITYK/MZrtG5xQOK03rAa+YW/
9Dpvvg3MsH2qI01as8FsBVLX3ldlux6pCmRUya7RIt9mkkccBXZB8fRtf+OIBB6S
fwvM4T8Mstk0leWW5BDZfE/C1v8RkqwsXL1+qAFFH9NcaWvQJaY5lpi8w3qOB04H
gptQIFrbbUVByqWUQym2yfsTDNZSaKHRoXaT5cITSUMSeBJqQp6dOaOEP5iW/TNi
m/pU78FGboEeW4FNemXL31yQ9aB98QT3KdRqz7+Xa8eAtWbPZr4z6WVwuXnPuOc4
qmKu/YFBNYEQeI6Ew7S1QMqpCnhnJ9FB817x933C/Gb8PnV3irvUWrO5/4wiH+Hf
OmmN4eprEv8i/frYjZrPhcV6OXlKR7/7LzzgABgQeTu2n3Bf1FrysBDMQp5NvVuL
ffOSULW+Pq2IxRm4NzrJxZOhGBFjAS/iuxunOCBHEcnhofxiz4aTNPXc8b8sMxCb
t4w/BTkJgYseKh0MpPgNIVJlvIvrEAL5LjSlfdzQ9pOMXSCH9ognz38kHysszvI0
8IGztsvshpob094FP3PmN90IyzlPB/D6osVUrJEmn3y4qgXrWoH8cinwtw50a8pT
2G90/RwEKRARo2x807RmxmsYP6PPm5XafPt+/CYdZuyWC7jRxWANYGbqkrdjonmb
pYbWYshZdtYM+KsbFREjLZqyIXBT8X+PcDIjqoNe/Hlr0jQ/AjhA96ZpB2ZMTYIy
6wbB9hZguXah3rmdzJyA60GZLr+BzBC1KwiTjSkULrAlYyb50a4G9x6P+I4StPf9
aXlPZJqCCd0NRhUfwV3gtz9FVdg4bviOJsTmnr+CziuEKBAGvkYm/N5mg4Z0da1e
Oa3x1lf1mZLDB4Wl0C1Sei5aGtwGSeCCQcaP7OdJg4xZlO+WnEFleTQ/pUSUj/Cq
dCwQPw0fndWE54qg0UYWXc6wYGgnkhjC3dCQ3RKBA5ubJV9LEnVdUhK/nWOfV42q
gXqEPO/+n7lTg3jgfFecGSLxSUORKQDqh7H05mSjWvbMqUXZVjmHr5xedRNvIp1n
rfoKORwZWlJ5nrI1rKx2NFR1tyiKWZB7WRCVzc2CXOirORKKHGJp7Yc3WeiJJrCy
VStZQj7CwOlRpIIDU+dW8uBuNCCqbkogCHx+K1br2LPWe691zoeKiLk9Ar4q4/H8
AqyMwYHrFQQRV2a59Oq6E+X7c/lbyf7x3bqrX7TNp3GNUw6BmsP7qH3yS111dVxq
4YLRscDGhKkgjt9Yma4EAjkgUkBZUjPxhQBT1NwPZhvfiFbGjj8rNKrNoIasRo68
EA16N+TRoVq1i38AZ/BZM3k47ZawjV88/xFj140G8Fnf6/Ech2Z142Fh725Z6jgZ
bNOwS+JC5DSZOwrXrUQ8ttiJjn1k0O/96wq6xJy20mQerrO37cqNkmhFx5pEltTG
kjFVMm909fetLVZiceHoy9B6gfDvW2hi0brndasRGQd3wQGRfwY8Pmy+MctZnc4w
sGjkCHj4leUVskngdmjA4BW+Htmy9UVCTExtqUlyXAFpiYjyl799L5qxkOnbJgQH
YNYSyH4T530Igl0uBDp5JAsRcaZCb4N5InDkwp3Q1ye6P3hmyTTdjoyO6S/39bGz
+J5Fn0DiQK+hTfyG1rFcRRRa+iB0V31pTvTrNB9jaBiGtSaRNzNDsz72otVPR4uA
x0TWJW2m98zrmL4e3OXSyRyQbhwuV+iUT0LnQz7LLUrrzVoXcb7ObYFXlxiGR2UG
TctFCyQ24WYM2P1opFQmhzTIBYw7W+M621kWbhVMOOjqjkq21f4mqhOM92ybvIgN
2F4PQ67517Oaf16dYdtyzel29lHgScKIu/jJSt34xN9gjSUfPz49JnMIiZQqL718
FqoNYiBsnpVCmOt7kPsefqNEP7ssewErP/2K3kOCMBQVU4+GB6yZVUBGn+vEYaWp
jk6m6ilYBlnxs/h5K9sXVumAQ29eLeAJEunSjg4Z3amSP9VM3RNp5+rmXYUX6ocl
YhXC4gNzGnreWK9qaDHsPV5zGfCr7OGqQR9CCmZvEunS7Ay50cKGQ9pgL7rHS4bo
8tR3Xt64r0/prlC4ubzrAZvcfFoON8Bry4QtbTlrIGh2lPyC5fsmUmzGRa9S9F7q
+8YqUMo8rvqQx5zGIuKuNM+SZvXFhg+Qq4Ui5MRt3OyDzCA7TmNAOS6bORiF/Skm
tdy46z368+0GI+3CTAClRQqmNQnM/fflroyXTigDWlVYsb8QGmq2TjarOxtQmWAf
9sS8ztuqHtGh4wTUrIubZQ1r1NwDyNTorMUcTwxbGYqzkltCxNENdTGibfMGkg9q
Qditk+BnryeAsWxtYz18wBYgh0Au0vHmocjffXxBVXju1zeyq16JlAHKC1WpOmp6
FhOAp5nokv412dawAS4zVKzsv7b8HIeMxWtz/W8qW6DjbhaIz7SWz87noFf5w1pc
fxxkv24tvVFd/UL5j8c27HhprHZxbjyLugNTmHOpY/Hpw6265neiSmRTa/KnkDjc
C2jpslFznfMHXbj81NXOBmj0eb9jUHwc7KEDblpRIgrVqGxu4UwB5X9ZHOAJkrqK
Jc+OVw0DslNNy0Usq14comPdLFOznKkZUoZ+iKZ4MPt1PpyVhjtPYCu6Urd/3OLC
9s7JQ65VEGCSrNzU5e8SXNXNNWNPa8fV7qIm8tylPO94T4r74bo/VxnAMBYsanX1
vyZ7CiO0RE8MoBicBee7+vpue8iSXGerr3+7U9udbM86y/rvbALT+ALIeYBFqEtL
sskTra40LvGK+QcxpH64UbWWHDmsmtRNR2LEceGYeueOYyAcuQ2IZ7SjIGSkfpNo
kcZ4cpbcnR3HW0TrT3xV+WxJttQW55H6jo4BpUk86bNoXdcbl+tnJP3YUtW4nkbK
gS2KHr7jQ2sMjql7L63GrVrGcCsKYuQdxxpYfECIBxJUBD8C/sMbc5+v54euVwff
QWJLo5DBSwSylqvdX+YDcIBfkO7OLOP8cEmqG1rg2v19FVXNkfDmurMGiClpBsQd
UF9c8TRyisXByWOiH0ounH/11YB6DSk9E0H3Ux2BghOD7KWfDa4BcjbfokWpiPZD
RG18nMG5BS024+aocYP5B2yuAWZVkTtvSS4N8kjDummouk1AamALdVTUbE3dp77h
rbu29Yd08dSGwadtaBRq+FmdgJz8IxpJj9Qc6O31Vuswas4F9gStoZmIKfL1CjnF
dY7sZBDj4/HxhhVFozGA0lE10ThTkyhD6qABJ9uKe6vPf9V+Wyev5khDOlZNiaY5
PCqjEwMkXmBKbqT5Y43CNVFN6/94bB7YuMEiJrvEqrytOXhWFCnkLMgZuSAWVTeI
OI1EyGC4UBlHP2+XPk5BAp+LcypsqhT1XHJ4+vsdLOYhkASii00Hz3x40lnbllFm
IjmY8+o98aSHI18/79qiRPMR8Tdkcq7fL9we3wxjDY2j+zNiFmqdd9Z/sSin04vs
m34v5dzbhyu89nXJGxiqHlzA7I+wPINJQ9BqWsShIKLsyuKK5skHdN3Rjio4z8ii
YerO8uOSVMm9pOxKVvqsZsC0YiLlblfqOZ1RWwkFwuqquXQfvDzG//KI+bSiHpa1
T270cIvloTv29WSoP/tSni/v11ulixPqy/ea0tvZpWpqmVPlds1ie8n1rS3NYW4X
alUm719wbUwZgcFtLcTSMh7yBpD3RiSMaX3oz6evzTnbxrVI6Qi4ILkNqiJiMqDI
uexqCPRSwRisSwlTu6dngVZU8GDe41TxIhm2fmnuvdPy7lkTjr1GAsgzW8/X/PF+
FtaYovTf+NbPSaeTYAJL6NI5BYahOwf2klDRLbbVXJl4xK1gzWb8VieHA/Kfracl
W9tdSAD/GJN/tUI+h8Hy4IX/OPPpnYouHwT0N8i95JdwBd/OQrZcRVLrHbRcpApX
5n7MbIFDiBwyTrva9Oaa6UtJ755RLl7f4TBPH9kwXcCOORzgIJabYzfu7nRofrMw
F4GOuTTbYUV8xVlhX+cvK7GV+OAZM6OOisA74LoNmCNGTORlYTT5PpYp/xBuCeB2
mjpogsdT/0icsUZqdJjatrNXYo/rmGrKzENtSX5x3U24MMm/2lI82zerGBjypTFF
7g0tlyDmwU83wJdXs54udQNwIg3uaxANL1DKDwHbSbpmkdruvuWgPHypVSr3gTRw
WzxnqC8ea3TzA0BcstWXoGklSjSmLmrreqAEIYZs3T1p8vWP0lVY6E9qAIw7pZCA
UgDiHa3FBi6aNf1ru02zf8ZESoq0JXw7V9l3al7yc/lejEQwk8kfUUx0OdwNoxje
OgvQhUk9K81BFYSjfFt5DO8hVN7HUmWoj0n+IgwFSQ47NAqmzFz142QQu+B/0tJf
yYyFW2QtUeG/Xsd7GkHC8mdJmHJU8ENKsNzxIjHsdS5okqolLz10VMCtrYfIWPDW
gBLvsQpwIzun5XmS8Q7K8RnjAOAKyCRCSHSYO38UT3T2SkWidqZiBcqlPh8N26+M
nct657NwO7/+pahM/Y+/FHAkxlrmLJspdxYXpu5w9oVewYmXPk3rmg4o6+O3u1nN
cyozeTk6JegmvMsadpuAG+I/9KuOZd918W+eJ7FP29uJV9p8FDaFAAQ2Uodzepoe
9cQ1Kt0dpbJa6vSzfTsEzc9Ip1BmOvgGH0cVFkaLotKj3uHV2xFcuNzGvoKIvBil
4bdwbtYOCtz6nGcl5EEXMkIFj6EQrRHHCWkvo6fxvfLbdxKIWVPgAtpSKuV8KsF0
ot35MoBQoFEZfGJF88DkitT+NiViXL9V/Embg9if6WlOAGgw6EA6tMebmgiU2q1i
e0bfxOGS5ib9EChe9zDIa2QqSVaaeomJpFusRSII12UN85xSSiZ+yY3StU/FyAKB
ZiE7CuMEbxiborSniSbSQAmWBHJoYe6RRmklZ7XRXjdpuWAWXzAgzLaoQgW/MXio
syZDRl36iBX4DveTkuj2nCAUlcWi/MvYjH2A/11Em1nnttZfPijz42KefZET+xos
L1mMXw/rS9zykfeL8QcwlmUeKsLHNEAMb4WNqqDIWUj/ivLZ1qgVpAs/Wh0OgNtJ
0OxzA9ZjuNAuf7nIO0W5nmV5qLOQ18yK2evVnkVn56k1+JC+V6JOf4tErhfA3UmD
9ALHx/6HPTQ4HHknI9kr8NybqMXS7zCwEMzZJyALVcMyrUYXz89EyzaYqpWWaN37
gr1pYJ5Rg+vTD96L0MxwMojAVR0B1E+wYoq76hIGbsBh+FNn2aLfTwK74EeWMBRR
pqY+F1DJ7XoRDaFrLW+aLq0LN822tr1wxRVU2EKariBBrs1fn0Mmu5snwUi6IH3C
M5yUL4YZm/rO0EvFQftYeoTxWNNe5XlwgBGMfk31VHibAtB3ZxrB1Jek+FFfshyH
E+qc28popbO1BpRwdsZT4VYo/FNY7m7Hmzl0OyC9bzc4FbY9gSZ11XaDgZrl9vZe
cAUKP3DCoMNXbgh8pqz+sy3+agR/JXu5oYec4/aTP4uOk0Ou7S3E0+arqhNgsVCU
tvC1raQEL+WCv0bb7b/47DYZCrWglVCdvuS9GNr4EGTkhgTd/d20pEegFYB0op/U
zu1bWqYbS/8TI8Ht7iUp2X3u/PbiFWSB3AXFyyDcFZBLoh05yk+OgCx8E8yGDqTp
mcztlDepG2ya6t37P2yUmD5rXYg4QhEYqaKHw2nMNgr5bxUfig53gXbLEvL0KaYG
huED0+bxGtDI5HxgLR+AnnLoM8CHbtXzW1na/1LMr+BCBMZluvAP8qdLZyKOjjdV
ojuWbEv1oM9SUhOHJj95JTICxgMfODxXcDMSzXLki7oRKkSrTIXINeteH1XzOd93
c/Nv5NSTGIaqP7b2P4rPNK2nDLIEwM4knvN7HwRI76tKfYm0lokDadvN9JlxH5z9
Zw2KgEoNobKVAKSSRbGVPXKdMAVaZQwtMsg7inHyryrBd1es+Ad4AOfmLYFm48Jn
LY4RV2Nx9M69/3s3aHvle3/YstWO4ys5yI2H3ZNI3ps5FkL42QecYMZJYt93NmwX
N2JTm+UW3NVcyx7I+6fJrS9IO+eSHPb+qFclY09l6jJf64VEbDDmmobZ7vJO2z/f
bHbNAs3g+76YvuvOAXATsecUPfKUapqOr5CwSrwqNlIdAjgqIq0VcpKgWdwaJymK
4HYAfHKK95zrnwtuUYqV2zcgwaN9YVF6su3+/UK3ZaKNtVwuqfA2JvAFVKJ6237D
Izprqu611DeuPRCqVi9Q5YCfD6nLPFvmf96CH60/QV5z6f603VkcrfwtqO0lUOPC
G9JDC4MabDtJJLF/DKMZAeEk6ZDi+xyVwvycF0r8lxlg0ZsNwNFGdLhXO7nqD4mE
OtdGY2XB0N9sSeYhSPCst00+V/4hZgFsQ8wCNoa0BxDCTsZIW+i8sH5mGvcGzqOD
qsB/8S8/fzDTn5zbcT0Zk7ptaRlQB5CgSuawBedtb8wRXluiXqFVzwDd5bQtOQRp
eE4DRRTOTNcJGW43DL48gTJbDjl1vHs6H0VqMr1cJhksAfS209sGi7iPP8gJCt7c
2lRcuuXwTXkcgLjjX5eSXYAb5iGwMlTOWYcA+JyvaaHUnBc8tJQ1G2FPs3aglL1c
IJi6qDNr3bIC0P5XVfU+KygSuQt4YC0e9ERkfRhExlK6TW12849ej/JsZyvoC+dZ
EGeEivJdsf372HGH+MXMjAc2MiipYIA5X0Y2WLNdNEvhA2UDZ5/OgUrvleRtEUG9
xG4Ufi4XvZXmN/YkgpGS7eZkM1zPSQAaoTWQXwrzBBOVar7Dgt0QPQ2GyTG6pKys
qCql3bpy2SE83Z49yYZp5C/hMhPOZwhXLNtZaNbaEmbgssTEzELm49OlWSYas2E2
fo9vdWbeDc5R/HraZ2Wkm7uVAbKxeRC/hV7zF4QhmLmNfy3s8ZzwdMIfZg2c6/fp
2f07JO3vrf1kziNm+oQjFfVV1JNcSq62dRRDp2UVYVPRAUPl+BMbhg3FWAID0FkO
3cbaWqfWqZvEMN/umr/cvPJf34rpUa7kYhoZDwCqgxfL2i+WNvFMGi0LcPZLUbdG
tj6/NDhHi7DDiVQAP/eakcj1KZhpTYISWpgo7HKECSVnH/p8vo/9upl7RkiYHeUO
I+V+JdVA1gHmRiMyMR6ml4l67fkwKQT+k0/MTPAjC48csLtU53cqx5cIKBCX6LLM
/1T70Si8x9yHju1rzIhkzyKdRwA2cPdGOVhOc/5kXRHWmXqeGX68mkReqZmZwyk5
IZrpA6LMcQZudiXWOwPp0efT4idBXpyscF/LcA4yCUTm7o+mZqYYaEGfdJ3tHX1b
1TqJ/nDmdEHGI7VlyvKOGv7O05Xrdi1TEhK1OxsUxXvgyVvbZcyaIBQIWk2rqBpY
cbaHpKhDqeVsbOoBySWL0iF6g0+5CR4ADpmshqI9/r0DQQ5cIJU7ScPsww1hXwql
q+tLO4g8fNWPY+IHLQUOgDFf+QJDwI2YV1KGa3lne+hGfOj1he4gQ527iMDpg0so
UX2nVcZ/5p/sEFaHcCtknj+DRakN2Gw4YoPBJCjzwTpMBvX9BR11XSE43BcHut4B
VURiO+n2IYeVwPuGVElDYMr5KtEZkvJj8KW0jI+kUo4HnJhQTPQ3oTkLjiC51Ynh
4FdJjmBFUIAG7i1tkACWsBG5K30gfvQvQUpQYOWenWUKEpFe84hmloPwfey+cTb7
cJEOEVZqtMp2ZVUzM0BHPnuCJN69tYHNLX2REOcdPII+3/5yBs6PkIdvCHoy55q/
pirrI7FtCqD/QmF4LhZ4H4utp7/5XOb20bulnQuMLdu7G9JM8odNHRrK/0HFAVxH
9cUmimrk8BotaBr83vw5bO6dJFGQ832WY3oOln7+oB5diqkCf3uP2RIlAvjFueqk
LMs2h7Pa5F7rzKwEpi8pyWJmwsbLdb1ePden9YkRueRB2nZwpvzuK1SmVNdaSlZM
zVFUD00xEg3FCa5nzEf5+MtdAMy64N9LVlmKSOdSuVbY6qN1/KiYFVXrtxiHnIVw
3/DQbpOfh/zlEBXDA+U6cB/+FphJgdWFJgLZKaHT87VNE7Jjl8IEs5iBiHbgdIDe
c93itNRLjd6bGo9JEslP2KWroRZaSSKGmc2V5xY3GX5DEGFCZZhE+r8hAvQmr1Lg
+WJeEKcqQOwkFi0CYaceJUKb3EO2P24NEy6kvaddZQm/TC7EmZcxU4/+VyDgw4t4
+X/feSDlmjzVPkqSHvv1TnCTGBfj1Bv/src6LsYQf/TvI+0Nh+BzK0M7DEQD5nVD
jRghh+nJd+Su9cntAtdfXJZ628+DW8gX1zLKZRZgfZzFjchxdBU/aNXahVB+O3H+
18uJts+IOlezwUhe5l8sG+hwoUXrjKxHmhV5s3sUJ33NogBHs4bFHEjgUjcmbAr8
uM0HRIIfugd5LFF/O1cSiR2uLGf5hexIpzF97r5MEZlsReABzc8LxqWjjNR/2cYz
2OSUxs/5hDOXaRFhew70rBR4P0N+6qZ4bPgPDO1bDn30PG1DpFc/Sdn0sizw3HXt
Qgg5CCKgI5O8eaOU9SkD+A71CNtXZI6kcbNlr4cDbwnAGpiozhj7CniIK29KLEo7
tKPDYSTV+tBnSPcl6syaIKMFEW85Ap8uziagGgO0VVaTHZRqYN+9thitRrbqtaqq
6rBC13/D3bx1FrAAW/4VUSitvB/oQEKNVxG8lXqWmCuqr7HXssg8GnzD9pIJtso9
avLmeS3wC4236q8kHdjklgFZTMUSne6yRft0FnruGH7bpaEUy7lZentCjEjXWfl9
oYjKN0qWbngOaDvNk9GergDyQUA81P7QQCo6kAtWFBQRIGioCtItBoJrV5EG+05Q
Cae2IUmH/lqR+nImr4lumHEF5aUDfJHcN5ALgKAQ3aocIHZYXmGPvj6LNqLPKVIb
+MH8rvU4CXjNPRefDjFJXbi1fTKHMtvfWqPy83D1D+wX3IJhVPFnIj7vmBYBI/S3
i/39WbymNizVQ9blkshheW1tYYrLJlVDp+G4sGg9U9mSjLqrv0JeO5Dl4fObKij/
2a33FKSetAz6S7IvCv1jbv1fn7qF+GbF+sNO2eWn2VC1QQgH1e3yiLx17oGqhIOq
wbA7OfhHXqMPQJ6WEvPtN/d/6RH3R4nptC10RRJ5aBWaI+NoB7XqA3PB0VeUIvbt
ZG5vchbRVKq/F1nlBiGWKwVdCs0O7RTrlvCBecytoexWPRoFNPdccyygcjXACqCb
4b7Ft0KQGNaSy0OrNbEdWOFwCrZh1ileTkl/StV4WmlKISyPsBs0n+3ag2aD4DFW
5Hf2R6YTefQ9JP4d7W6v3rDg84J/H+Cl3Yk+exU15n5ASn76ecTSk7i+Bt6gV4pr
/fpD8wbVXhA89EPvH4C/5YsZKPDw1l6rFHGuQvyZo1xJYcyk3loQygmJAuz0q2mF
cgQSmKxl1Tv0vr/C+lsRcjNPDY7j+sgXtF49pT+0IiG+SD3gQHRKCtXlL3qvuRXq
yLsCCa6v8s/oiqNQEpV4hkvTJZfblU1FAnpyIIpFFLXaJdqfNXDuKLQLv+aLDYvP
o4oMXJmLqguWzDv5ygyOTg/n4vCyAkzMf1e8eMm3peNyxgstGPH6FZN7lwMrQA4z
pzwZL6EEB9Lygazbgnx9m2Uv0+vihB8cHU/ZEzPR+fsYD7cOPHD/8jeZQT3UDd6K
N76YNl7jrZ3MwEGRH/ELj8WvBj332QlfI1fgd+TSZkKtZmBOhrJX0imB8lig9hFh
RSEMhD8ZEoX5tB8rhFlaDAFJK8wQuevtMOJyuNWoY7DROv+9rJY35ACcYJN08vZX
jeS9ql8syDbzgZ+/X82YXsYya38UyyT4o2ELcNfZjYKSmXs9HN2w71bEYktvztxT
TqrP3c6cRUK6q7ju/qosdEh6oxtUxltLFkTjUza91HxJ6hDSjl/LnlLEZY25Qz0X
Cts70Gdz4JcrIePiaLo2TLt8x74Q8mBml+tjcPy+PKZP3q24M0qkQFX2GL9QStmL
nd22ttsrEfmyxUK5CU6zPBBmjN9k1ES0/K/4zY9kelmyNwdTwREPkQFguzRzzmMY
juXB9iIDCRZa5mLZbASkcE7ZJoWBx/Vh8XztRcdFL9BFwZ9kll3GoaXH4wacGnXD
Na/EUgmGPoxM1VhGLNnidcemQMTDCFgonBTcsPMd5j8jvKMM+LcMXcmtdcIujpRu
jC9tJyfBW6I7RSW7GDMjRB8GNq47Vxc39aYiamo/u4+q3rfmiXkPOgYvvQxrQfHO
Gs/sqkLXaA6MjFuJsYjizooMkpcb+LZH67w+MBV8a7u0G9k/JOQEcuj6W5NSYgA9
nfqpdJjE/aBaT54lzVc7dzkt7+iDQgNTLa0GorIm9V0bLctnc4RfWKNjMBB4idz4
1DgTjiX+jNj1QES3jPdMtFqwxTs8+9KeLOjg9WJilEU59bRrmzq+P2MFHld2iBhP
M9V0N5yf/mzeNnQzEhzaFHbTsAYq2ieQy9hhvNNVbSgE8ANfEeWGtmd9ltxp5w7h
VOsJvSWGGvTzId69FAZRO9IhxIY/P0jSy27D1torKel4KctXNwm58HJ4gbKNIEaJ
eKFkryjGpB+mBxz4IUhu+vdDefXp9cG2yoqErbqa14E6akOkYVv/k80D1lAS3wYR
UQzOadJTlD7hYjJ5+eU1sW5qiFmMzSdIAPwQz6XrlaTa32p59FQxUyFeXfAL0mup
OGGHUxzjKSK7tkDzFnw1XzdK+WDpTSYNparD8IYud/SrjgW8MLDXRFH5mI7Hb4fb
MuUFYP97k90eadzTJhBPHNQ56tgFWiNSLGnq/D+mMldrC0asrGBr6DgBLJ7SruHm
4OH0lGcO0l9EaXDH6esLk+tiVT/2Ys3IDzgczit/lbrh9nhkBdt7K3DsS9PXb/G+
xzMmdF5vgHmAJCGw0JE32KXq9MJvdeoWgiZMEZcB2RWSAsdSDKSeGIKHk6h5kALR
nc+WpLH93/LieeyAn4vrU1FCk78S+sXFQGVrCCXKkG0PxEuqktOsWurTtJcCFoog
r/50/66gPnE+sAEqThofzscZAhxahMrJJ9yStfG2j0VgBYtfnWPJRJPWemeLVeUF
l5Ui2EAY2Ywz2USwW6GWR7qExJgd3aKlHqoXQIKQ6YOlHCZJqtLA4AT2cugKLZ8B
MnkIra51+AN6PxZXmR3Tbubob/u8LiOkbKLv5LJNT1E6y+r4Dug4kwwiQIq75Nvt
3Qf29uiGsNAznE/Ed1Oj5PwOys4KLkKuVBhPloDfnSUkya0hrgiaG6Wu8REVtbKa
hVfZbTumwcItkfyF5PIB9UlSRJQGJxuwJhcyulFdxZaeX0pxxndMT8ccRl2onWQ8
kyytBQF+QRn19/Lk0T11QUIsz46D9v7Ps0Qr/cmU+pWd2mEtJEt4CC3avbLdgWzI
uGjfsldbYrpR5R4uXjndDTt3P+gY7pn2UGTcBNEsSsQ9QYoziASaPM2PtrLIx/L1
YKGZPfDXnb/YLzZm7JDAbvqT6GVlIQLYeZbSOjHu07LnS09YKVCNR0lWN0dpF3Ii
roNexrabWI0MS6ZfG3LH8GaobDiYA86JbzcFOnwQ2ogt2RTKaIM30ONxLxlmL2nb
I1OtBwViqEfOHuKjKRCnkZUx4FPPPdfIbF/npdT/sAvuk0lwXlKMSt+3v2jUsZ3x
iQXOeZ5IqbTWff10G9HDea5nynz377QWmymAALtpZaygcj6ZneL4R1BtZ6n4Yn/4
Iqg7O8hciu7edguR0xvQZexKxBCMjdZhQiw2XmQUtabwF1pNF1WpOvReeJAWNcfD
shnowos7XpLdrrL1tRR90Z7IsMeslFqW+Dcx1uMVUdkdcjj0E4FuKhlKouEFc6+y
zrOhApsp1OMMbpG3qCgDcw4TY3urdLAEFPivVZSCudpCf5prc1eOFHnBL5SaPfUq
W/g/1n2fKSvUNaAYeo9mHH6kcryvbcDf5JbuWRA9da8VD2n9QB2JX5Q0rWQXvgXG
X5D7c0KUdRfQTR5IhULeUsd/5KA9Kz+h2Rg03ODtzCRQO5jXh9U3fvxK+BfbGmRG
uX16GWyfdYadMNCw9pctoRzZyFCrIRZfxmZTROq0DoWgYEM5A4IxpVaIxoku9AdI
EsPexPNOATHmd5rzySemp6Rj70XUrgm8kOjpeHY0eWMjJMfL1GPuPk78NHs0DgOi
QjbuBfO8nnyhJfgBkIYivkp57KMd9615LW9Qgx+RYB7iiDJcZWy+/KplQ8x9NZ/R
SPzwyzh0dvnRUoNXbMDHrjOAKXZ2siAIKnBxBLa90nLirdSThh7o5X8P1+cDTnIS
7tvNLk9uJZnmt6ihaHc85ENKi3XxFdhIGBKsPO1Cb7f1TWwmciVssAcRnF3u+AUY
m+V9l8oHuLxkBodXqXwWrzrsLQBTzI/DsXMbFQhYwVWgbkKhq32QMQ/EAnW6G67J
MpzdzxILvLK6CdJM8JSJ6ccSQsMaCQnnVRuioVOhO8XCQb7+ZxM7xF9ZJXzFbsXF
wMy829XcTXCxAO21/jts/H3Jkg1OY5yQGlR22oaUJrAt0Izet3io0wS9mtEwx9T/
qnFHzv8hD0LDNTgNveZd1N7c+aGE7lEjXWNF1c7xri8sxyRuaAMbMr3KINY6PTyn
I8gzgOiXqoNSwLky7LB9yhy+wFPXBgpMKkHET/GSlP+NJtozELqoW36tdYI21rxx
jDPN1JRSPqDtK08/6GFUaBs1QHBawL0Ee6YMpr/AF7umlAjohgEKvhyIJ6WCW22j
RTqaBFFYRTDC/MWk6yIAA7RXBfstAYipFwGq0lWec7IUcmIaekZ9lhXBzxHoqYIA
NYP0UkgG2dpeFv+kflugbrGQ39KuScC2A7Wna8CVirHxLR0P1phZFSSNA8/KASGQ
vUSnk6ze6EcXgSbWO8+x2824l/Yeo17h7/tvsVc1zfN1rHFeT/Dr9quz5053nSYN
/oGWcFm5gbX/hK89bPW6JDftKqHtMfzAcxPHxn2xtk4NJBcykbYdoYw6PbDx6I7Z
h1hxMcVTI0j3gjYjTISNPFJtYUF6TTH5LYIfrn59dVgHKjVmwIWtIudxeKYgP4KC
houySHTMmLMx0z5M9/zRmVQPxFLwSs6gIZTJna6fAltjq/i0qKH4sMPH2QkvIDsl
DYkYLLcp0RS07KYcM62ouVLoqwQoTvnx1V8BeGBP0z7RMvGTYo1GlyihvMZWEDn8
UBUxv40mpDs2eyHzX6l4cfyBFlpJFmdrUQM7df7X06OLMRDER6KyHalNDBeOuCpc
prbkCEfKf/oYbA/QsjK+YIq4guHdsZMlMM208ny8IGQ9+e2l7m3MvjxTJs8wSEiB
98xKjIm+RSlad11fgPwNsRzijWem1wgWlI+rsNBvD9GRTRYVZ/lSbqUNb2BiD9Hs
ittc1t50uKpSVSA9PZmlB/IvsMFQBwsDKOyE2Uai2s8Z07N86dhX8T7Jm1J/pFeZ
X6AmMtI+Wzcy11Ejo1UkIg+PpcsfaeQzvGY2y/icJq8gQRSM+WWfG+L7TMOTm3Tc
fkINocf2lSaCjvZ9HKLKb5VlcVwBscRUpkyUbKjMnDNtZ/7ID+YFwzCP7sV94Tgr
0120r13GZ9HkaAHfdoaj6ftpSszTPJkbFTgFQyMMuhKov1J/iVMP/GKE1T3PeI3e
Hp+CgvcabMUeymR56vS9ezRkZB4i4bpdhfyDv043JkUeo/3XyBuQoD2YkZD3uHSO
Tvd0rrrgWCEsYvUmRaKnf9QkzSrebE0ebehUnxiLKdsEFO/P+1cmeoM9m/ri1jbF
yx9qGAhoZ/uYkAwlxgtM42j7b61B/CGSv7PupuIrN5Igj6HF2jxv5Wl5+9DhF6f7
apzI3t7ZdY3r5vg3X/HbK9RkfMbk/KQZKaAVmTLiEGhEVZx0vzFfo/UHYbm2ngv9
PNGGLYb6fjj4kgUONSO4HPCGfVSy7T2NU5t8DsxUMifWax/lLeLwcQ4jff3rnupR
/6lx6yzy7URt4ztoa6eHmM+Es0Pb8t55zJelb3MMzXJKVwu3Gfk6iIGrKx4aiDcA
t6UFdiQQAhe4J9wPdTlHgnPRZecwpzkCj+oc3GU+s3aHw+oVjQ2bymXcgrF6miDY
nJORvCUUI8LAl7+iOUfkAxH6PPeS2RIxrwGvoi3QBvoJpydHRhJvMgP+e+vZjA5b
dWdC69x3A7qQujm9QkmekxMDKWpoGC5wqy4JEXuGFQLFl7klA0gvDfuOPCU4gIgC
bZqmMS4n0HjKM+vTPB7k5f87ExVtSnW40NiMdWrHHv8v2fLTZeGkdZnZDv4Fp5aN
mv40nb/VOL0PU1WUT2uwyZeWKHKb0Q+03DTF0moi4NDes97mA6/1VIVUYwP35sQj
MfoVDS+vntBQmNzajWHE6QfH9Ng8JpuwEdq2Hd3MAwLbX7uZupC0QQp35Fn7u+oj
aoKU/OLPpv+gaSdMWneq/hRIXzSQR/bGtJZctrlv/EtE5uGjN8PGYAJXEZ98qJpm
gciaF7hvmBwqUGHi8CnIl/tuUden5Lx+HR1L4++8t4n/y0ppJI8F7djV13NcPUWi
lXr5ffSAJsCGY/Bgkb9dMmwYnbISBTMXMNbHO+Z/B4vIYRmccrtlFUDKVv3/p6CU
9w48myRjbEHz4ixKTQG1cLPtG4noGcCCzqtPZl4lk9GwgrpPMG8J7+h82auxNxcR
zadvRe5YlLvypUvWZiA1KLut0XYL8u6d2jL/yeQTF6xrw8V1INkofZkDZp+XWTa9
+zOfLb4JCXEgINGKavkBnIC836e2R6HIztl6bqkiGUqQ1/s+rJoCw191NOsERMzp
XyN7JctgBeqLdZA1ZyS9I4tqJPrVRwqoN11+uwayLrDgdCYFH+qOIqNsz4maoz44
o1Ae4lHg/l9VuwDCGh9s5XqGPzLAM/jvrl958Gto6n3FKW2uc++4eRt3/ELo0VvA
Cl+7ckdYej86hJSRNDTOpZY25XbwH44sUfboRvq+iS6kDnVAz4lFnb86lBwbT0Op
FKi2msQ/F/6SggGvqsLL4z2kw8U64Adi7srmdImdAmrYP1kyC803z9bl1o4G+4qx
7JK/J96QrbDs8P3AanpmGjC4L+TrFR0DhL9ucp4KyuRBt0gIvrbk4kJmX1hleWW5
AcMHadTAaRIC82K3T2cN5YhP13ve5/gWCVbwAoahiI2RxEF3Jzfi1+IJrjguCqpm
Qs77QLNrV609IGX5ZRB97z0vr2OzDjKWNaODKyIuGH+iW7yA63OfUr2vps6yeR9g
g3wq/Dzk4fA3XI0/nzm0Vl/u3c5L4lhDKoLs5ZcDTnndJBPZ++AjCWjsy6JZT9Du
1ZZ6JcWz7OPTiAkilhqKYYYc+DTmYsoCB16IKU8oh4mXIPH/hwwBfeMdUhY1VPE6
5l9zc6HbQnXCjKT3RnA2SuAUvZDOJ4J14s/9R2r8+WXIsD1otYXe3sZ59EhwN3Bx
ZTJiMs95grQ2teFgQhKTTsN/Xrod+/JQiIMi/5Nk4Jg0EU5evi0BhowiX4GZoYiD
XX86jCEAOIE/ZA16S8GwwM7/PVhY6uRxTI5Od9ycCBs+ecIs7T7fu3eX5ye/5Y7q
/Y+ZTy4ueSfDpA2XgZ9oGQZriN0ExCQH/tenwNTK3da1JRVPebUAjRHlzIKO5Cvv
xmLHcTVUnaOeC80tHVUotrfCsZj7kCdt5vpDKnm0pxjA44LTTZUV99ne5mcJS+Vh
GcEh96bSjB/fvEwedNelnojXl5+id4TWiyU+IGQZAhq8Y+wqqaBoAkk3/coioOni
FN7tan6LzK9BsGH+C2w6EAsQoR5lsCUso4K8U8KyPpac5NOTM1Sa8Cw79yVZRjVM
3pj5rsS27vGK35+L/ml6nrxTkcdNlEhWzkHlCNF5ld8Q0Fln3XZv14Dl0Dlneflf
d44FDWA2iIr69IMWJ5MZ+hPy8XGVfNgcoSIezf4PqYhAevMhmf1IHkG+NeqzW4NU
YIuvnSIsL1TBhOslojYDWiO326XXYrGz9LfOMlgAZ0dCECQ1v6UsA7s3DEr9evjf
X/EXgJLRIQnml2GV4GJPRGRXLoQ0rpjED+mMtpOCIM9Eb7LQK8uBfx8NcLNi7XNf
fIZu2ll04IcUuu3kq9sb7fX6g1NRhg3mjsoM0koIVl38Dy5od2YzVVOHjuhG1nJa
elClMDnIkSklwzd6Z9LwffKd2Y7++pnRSvCxc6TIP02DN2kRqySChED3ELpsK+k+
hFYMDkSHRgrpsBOpbw2/feN05C6z3lxh/DoAMlV0bl18CAvFab1EsWvelAOsylsU
h+pSkdiWszlrBtEqvP+1pR07JT3cQol7Z55wYDL4bEwStLaHUnke2oiuFkNHVkod
qpi6Vg8+/gmG5VKkja4y96xd5eb0ZBGS4HVvVCaszQpvuExlpti7qcyn0PB5YBvt
WrQvo/qBbQLvMeoJ4qnWTep9oKUZWjT3ddBJ+6hJqy6QKWH/66Wax4WS1YAPestF
MkYo/IkOP25IAE6OmeFoh0jLNEiQZ0W6t3OdsLcMmyNJSSLVH2sB1Do8ZyWoARPK
6OKaarVED75X2KnLLQiKpVn8P2Oge7sD5VoVyhsvXr68DGPTFWmebAASC0ivylTf
t22MNugMxDGaqrDlfNPeAIMskt96IXz/UmDYjEPZ2fdrVk8jy36hZU17K7Xjv0/z
sVl9uBGewtQJ5b1ns/lkjcH1wVnZCPWobpR/twb28LcISG5cgWFUz/i76hdjrQQ5
J/ODArJcch1IVfHbx8fmQY+FDS1bhOw0JEM9Bkqu9U+QB4y9lu+yqn494PZ0G9qh
fB8//inJYTZyiwfEMWU9EkDsSwN97Ky0fSUKHPzZfNA1fiOCZePUJn1U9znp+3D0
E3mDdi3g2r5FqklSbErWCOjL9zfYG9d5p4asse8Efzd6XauLkSK37sPq9RNI75Vt
QQGO51CiAqpbTGPYm/2W1ujMrQmlQQ2mELLAAoDYEWmbq0kWCs/iVcMd9a6lAsiV
FfFbLNf+DeJaC75WSOHmLG51JLQor2J/E1QMfOVwCxC6pKRYWd8ymGwmnCzo6qK5
Y0kJKllXJORu+uUh6EyIUH27UIDDRFB1/BpKhGnNzEali8F2h8hYWQEQ3QtjwfG2
2Ls3cCpHBzRUPxlNpBlgNbh7FjWihvGA7guG7qw6MRHiZJzPoW4Bj1kB9DJdTX+D
INZEznRisyYMg3Xv3WR/NUD1UCINyvK8MQGZ1ZwbVXYVzy/C4M5xMV0RxuwGza4G
w0oiGYY66XQP3uKHLQtgFktHQW8XEIT2tD5/plRqq5MDZL5bwswxm3XAIyoGIz8N
1Zib4Vo1r8TMhzve0qQBJaiXkA1a4dwJt37MM8O1BRDCQ/RnAtNcJJLdHr754oyD
KfV2MqwnM1fl9yllXcHzcpn6rVKzThNkrdCMYMJv2BloV5ELLRnzNY+Pa1MCyeXE
lmFcJWZNAp7SzXqAfkpW1iZhp/f2EJh4E0rxBUXitwq8RfdSZVcWjPJRGBeM/8+W
S8oAso7KrY5DhUZzGmM6d+uoe5Q0i2Prc2074RlUaapPKpQPvFApOVUNzqxDUrVF
UpKzFAr3nilTSd0/JQkkw7YR4ANHCxGRoAtxX1DnZPZOhV5dILPmqD0mtFye5Gb6
EMjlzvDp4v42HxIVbQ8NptZo086ouZ0i2PBNNHtbsB7PTOgXF5MQ8r7ZGAMSiy8w
JfaVzKCgJvjEzC4FrY9gNKj7PfE/RoeqSGIQ3YuB2Kq+8Px5CYPAi3+6JpNIOQDM
GDls4Q63TfGQmTQk4Ymo0/PJw6GG2y4T38FS4a+kxHUqUSXMH1Ka62O0ztApLbXK
W8Fh+KFYrmfUV3Rj3/0wkhWHIY5O/Jx3IeHiG2WCj8kL4NdOzd1v5iXHAzQrkvwo
+FTG4BYnHZrbX2NYoNLqCYrM7KlPCc/DAYwDXjG0lTCOZ0J0AYcr+b11fLD/ovTM
tfY91vEmCs4E2DknIFk4sK+nZS1c/sY1XbgZWyCI8TuxAvjd+hnLGTgr33xMl83m
9aCEu/Dg4vf0ExH1wust/at3vt6kIklu7Ny7vdEr69NIJrny4ACHf9mDsz8lm1ey
457JyzpHEw068rjn6b8kN2bx9KB0mZSpyKUWGyjsVO6bKLXoQcx4EbH3CkRB0gMS
ZmvGT2C0dQzfJTK601/hofUKx2zSp5VyOQ553O5aSSmqzl04MpCMkV6Sh7TFlNPc
oUROnxEFXa3t9wx3NiJrpM4VUk24WVVHUDhNey/M3RPStAuIDgdFJks9ievX8rJU
7pRrUl8mG1BuiiH6diaCUNRe3BzEE+xNlpAAJklVukvm/fKeTR62Hl4gQJr0jEI/
dWbX91IiujNEMSKEFtsvkkqYbrHa9GuXbgqegkbh3er3MduRZ10aAWEqDUymqnyS
D7G8DoxkRa71Md4dczpIzo9BJfCIFB/ulp8ymhveUQ27rOexmbTXH6PZh4V/rB0q
VXeNYk8DlDOozWQ23mbDNaYOUC0xUWp3bIR1ShGCDmLkAd9IQTmHlG+BDc9mXLuF
BWHxxPPqmq8Z0sAYSJ3xkIMxTm9VENrUfvAcVa20lUpxsx0gQYscgwBsGMFTeZJD
UaSm3zs/8uEhsqaDpgPD4gs8SPgjeoRp6qx82SC9AZJDbCe15JRBxwRYtPQgwXqP
/RexAl8h1/2QwVZRtBKJOFaW9qiqjG7+SP2l2HOx5g3TZp2eTK32BF6q0DYLoSSH
cdRxHDbo8RZh6hkJcK5tmT9NYZE/eeTzVyFlTeqctNj/SreUPQF/iGY4LHJGKuog
Fh8issMqXEc9DehysWrQSeMSnelzmr+zdYAJvPomO2lse7nRpL96YlWE+NHUJ7ri
CqzAQnPTjFZPUeb3z3Xho2DwR+7gYYy7Y+QlN5n0nGROdrRdVHRWH46rb8Iu67Gc
oP9QA1Yv1eVNy+LuaROyYFC3enq8NCBaGOvGbzoMjEqNk+nmBCa2sM/SzGbqerL7
DNc1UURmYrmAdpSWrDFF0GqHAt1ABtnGfnC84HJVrRu0BgT/Tvuy6GLnPkVNC530
5Hjl86YNAaaVgQp8tWgkom/T89Ec0jNTJNH4Uryhb+FPRAYJqvU41pyRdUZYh5fJ
zaC00BeaQuITAvD3Cj6huhNabPskIbxhmjSlSZFIcOm967SFqv3oYhY45bUCwsC+
YvhrGaIXWB/R0MN/7mlDTwsCB/D/ZjzU5L7ONm8q1FOtHyqxrTVUYu0cULYC20y+
IDw+QfyPukCswZq1rBGe893+OCgvILPBEkKvopEhnZqUYDgVoWhOyk8tOJ1nivHN
xdo3RzIX3CWyf2dntS1uOfAjBNif+evqx6iKIc2YT0sUaEtQg6Fj8R2qoFKxfWP7
I3jGt6b0feRGBzzcEvMonuqRfUO3CqyvTLLlZyJCqLDsFtn8MRvWOLt0jfoeqMwh
oS6WXxYM0/BpBK7UghZrcdeIc/jftsqEUc2UxwW9htMYZeDQETErB7mVWMj/Ab73
SOst5vYoaTEie82FexzpGS60ZO8Fg6O5IMhRW9Q7ZhliwwMB/DL9WoSRD0+JaoMw
F/fuJIwSYXsH6BEiSnci1UXsmxWd5KEHPFl5OpAyy9WZoOHMR5x08lHpABSB/aq+
EDg6oN7AfrY1O+1g+YItIh7qkronMJa/Kbkm/acUcLDKjyHNnYsnrpXtGrYe+6K+
mpyiiFyo38IuGsULwv9DEPwGyiupnBBNRs1SO4Yy1qq0zK5iuv0ykOQlF7NW76k+
Jfe/dFCv8lap5R88lSSobr76Gmcht0simbauaiJLWEiqhx9P/NP08MkR4PMLsAec
3lMWlLo0jFBGm/fZFih6o9vdLCV9DfWsJ33nP0L6MgVpcDAZUCCw99cuApoGseFi
EuBRGCJiFaHnYQrl/Xw3lijRcNcRqQDLhFkSa7dTfOY6GdbCDH2rx6KQbLXMNK9P
y+VrAGB6miKdYPBiC3EmhJqYTS5O0Z0VcL/F319hiizWGderd1a84UhDDwzEn+Yl
5ZSHmX2G111VxGuAuGoTS3vSJn7UCFQGzUJyg739KToTaB/dTfsXjOarFJncx2sR
08Q7fis89dYjNweoupnwLLAeR9YMM0kk17XQFITVIGdtey1kUItPz4Eb9BLDkmyS
xzS/YDANwO2N6vNw3m4LBtrPXkuxwu97cWAIKbLy1NXRKWAvmaL9KlcgHnHQvVux
rXIjQ2XzmNlQzD1esile+ouMwkmIn/op5KlqHpMn22yVKQIdEjy9dluawC3rmPJo
Ir05/thDOMPTnDIF7Nef8X/wwWszsqimbMKN9LCsKU5o7+DB4J+pYdnlKfgiiIHl
fsscM+72AznCOfQ6/WI03GR2d+ubPfjkKTlOktygpwcAavp5pICB341/JdkC/emp
XKBFXFS07gGhxllHqdS4TflYq5RKlXLGNDjXInfochzWxptaQC69Pabe1TUUy8oP
4AWRZtupnvvDUH15s1V12j3pl++SJsHWA3e3QdMPsepUM1kw74Fu+f1sGsprWY31
Wf4rhR4UETD+8u5VOXuWy2oR5/ICpAV06shxs+wW3TzPr/ifbNeQS+dN+Bum1//f
sNobM5Ox5uTG4Abv3xk/IxdSAWtTdF9XoIvbO7HQfBqUBZLaiIqa/AENrV9Sl5Oh
D9OPQWN00lG/KsKn4+IHCbQfHs1kQe2wRVt/WmaBY8M0xQCVoUAXyKlOYcUHcUA9
zKgU/5OuF9o7FHx0qznx8dguVqT/Mm9Gxzt/V3DrA8EFvkxARBNZ8SCjXsUJXngb
FYN2nC9DG6NKn4wbFrMbDhtFOfbAZSWcY3fffqs1FuL13MJHCcoHpJ03YWZdSePR
GiWfohFLjByECEhtqal9QwqX4A+GKTpt1bjKQrWLrfoLRj9jnd2FWp0EDAargJqI
s6oYegR8dNvhptLHE66Yuo+ytF31WCCfAfekKwfaKhekpks9rgJ1eBwLJ5l21thI
hurpKhWL1Gq/r3d+N6XDeQHEMvlmNTMfAK5HEsAip+tRf9ZLzd0okT15Gd1y8xZC
cjXAiRIqzLw3gzTGPFCgmlbN0zngTYO4RpGAUubAJzH5Q1X55AWxSnweii677XAx
hCCwEnrBN6l1ge/rrtFUgYbBCzdy4ylSH5Mvat/hyEt2GYLX2aMUYuYP0QRHQrW9
g0JfgUyyJbvaN7RHelF/24DtREoIDKGOtr0wgyYhcHx2JacUyvcPZX8+fnzbsu5+
F+b9mWFwau/UHGOWHoFwe4Fy5qiKsskMnGn1BRgo09/HxxSwQjwIJLKwOS61KIxr
FwNqV9RxFlOmozQpOhm4AJ72z3/Wk5tWaZcGtBVeGNJc4yKJrRkDvSXU85Du925J
Ee+6wdsQYIzBbyLnCbb7Jt6P6lA9mf6CwTWr4a9/x2Ce8dZIOT7ipAi2TJeQoDyA
YNgOEUnfWiYNGKf8a0PMeAIYnWiMf9OMBb49s75Gk0fewtpY+gRyKgoeH5bjYQ4d
grcWQRUZWpfKOvQDflX8vY+pOgXz7Nn1vXuv6rs5l6ossniWZ427EGlY8Uqx2055
C/eXtJ1VUQIwSbgWWT25nLIlSu2dd39y9HQGcxbXCLbI5LTJ+sgSIv30vFRIxJZf
2aZAq7MoQR5lMFHlSeieRREWuHSCSgajI+6UhrovgQVniZ96upUoshdSYYiZnJ9D
NFrmG8AbJ55qsLC6EfEXQPIWLXpHDfkJ0M0tPV/KvYpGXYstTT5xqdwhRSzV0q8E
lAyAIQY6THYmsfSIxCyAj8zTjVLSRO/Pmt+eurajQxqmXIt5Ua/onrjaS+Wg1ju7
cEfpfyrM6pspUuJANewhgUALTjTld4jGICMwWsD1RD4Dss0UYJK3skOPGOyNwHgj
+e2kgCCmrmOKfV7bHqacTvRWlcMTTyBGhS6PrU5gbA4HBOIP3+sgiEv9NLeV3Yht
7RN9yBSaxGwG3PEqMfUEoLQhLa1Jydx2tcsg/xJAHwpf6qgt0LnI0NpTrVprSgfg
8pl4MLiP257pkwL20NUVFHp9ZbIMe9KoYuDhNgwGnUjvfLJxZBxRVEt7ts1IjuiU
BNvY60MQCYDNoKnWUY/ssKAgw8zKR/BTYAdw0wPVsHnS4J+X2pT4dUEXHkMsSC4M
K43lUoHJFiclcM3AQzoFOD2GqOvT/SFIeTbLzCqbqhX8OM+AHpzsB6EommMaO95n
qYGvfrz/Z/pnzimCEWLr3+04xsEAptcazv9hkB7LlI3wO/VphkrPMm6P+NHD6kZV
2ewKHTo+CI+lYyRjR9XSmGA8DoKfzUxAj/huyEV63QSg2ygWObQgHetT9oSNZBQ2
Von9E+wuFUTWqdx1zd/DxsGr4XVK4MZTyIXFGepVpFnh/ve0Rr/6uZ4pMAumLuNH
e6Py1Ljq6TadA6KYxx/XlhaSEidME1qxc0Y/+Ra95zKdxvigl5mCOBt3TOn69hOw
GehzO5Yj4wsV3qhI5557pmLVtJfgDKvJ47Nk8GI9XnPg4Y24nMNeXTfZF/IX61sE
fsEJ+fGez9ay4sX1cxjcPTsJX+4mIub63VIjY2AnwEDPmMliilL+0MkS0xZ2zX7/
463eobI7x4EDZIi/TEfOG1UCxUK+YYwECCiYz0qPrqGEah8rw/wd67CM7BBEKTen
hrHErkt54QKMks0ZxLBuqW3uCrD92m1NW7bDqRPM5ukwwtn8WZL2jSSDxFRxC3fk
gsd90oZ1o2JmiM5iOQrCR4dUtvxZwSYtZ2s+1XembHPnfpNrUkfF2Lq3eHOK1vQi
US2KyBbGgghEN/MYW6TbLZdouvk471B1RIM/ZmWB/ntEoNM7OPRw3wwld2Tz0hAo
L/OYW6E/4eblfzGSBNdGClMEnXkzRslxFnWf/aVveMm0J7mpVEyqd57deTfIxU3a
bmj42WeOgeuQkPDWIX8w9J5g4fgK8vnDi3RykiC6kEB1oUGsUem7WPMT7TAOFMFh
I8OE1sQgDg0islE23d6Znt0EW9IAuUCUHfrG9FhWXUBGlBqzudGCxPMlehT9E+XF
c75LqIRangyaiQj9VEFTiJEABsE2LAdEv6AdiC8sGkEH5Bq3kVniRCD1LKw3wD0O
PUI6+WAYd/LLxAhJg3Lr+7F555+ykH2ryR7iklO3Vm1JiTo+5xv4gllthyUX5tzG
DqsXFH/p8RnplsqS3h/6G7VlCCZwpYAAyuEYwcsGPvDC1mcKDnJZoFgIUHr3Pnul
NaHA0qe+US40U9jcD0HdiROgCZ7T7vOwZMQ8OaNz4/L2PUHFpEBeZ08VFz3+qTfH
BbOUDJGrQ6q9sAcMuNvRMhbD87oVrWf7iuC1AVI28hpoMWI8Kizj1MWu/2MkdiCK
LTEPWGltTrAEs7XrrwSClgL5Ryv5G4ddKJI6Pdz2/8GAKX7AMsvUxLmAwgoDrzZz
wdufeMII1Khu9YXT4j764ZnlQUjJS+bxMH0JQ5acKgIee1y1gWadduBeP+wtFQe/
CMT1s84oeRtJYr2jdjFcD/2UdYhbFEEvFa/MfRmiQ6fXBH5+vLRk954tllNXciCv
/xuiYgyV0mRFKx+f2qn2oUT9QEZL3w7757Qmmyx61bJRT9LuPii7y0edgcvDMdF2
0yNOmvZypIi7MoDuVA9h8vcZ5c+1Baegk76x2iB6To/ymoHydc+o/8wQ2nlTneHL
SCJhCWiyAxpVjNmFO+tsUlNf9BxAQCSTBv23VrCgCpj2628iAIo29loUKG+29F/O
6q0OYlrmFsPrpc/pCOUxftGhwwv9QCUAOqzzOqCbQBvhj5eLoJLl9/vdULiB9LfU
+Ex7RTAXpuwIVa/6cQJOjYUo0s7h07Op6aHejG3tnRv3dK1QC5gxQO3lNwaiuVjN
PdNFy2rncNc6tz7MarmBkLb7B9vpio4+SiSaX6SP+cAeO9YZCKiC2WaH8Q2WWNbZ
RqNrBvYb27F5MeuHdlZJDsNM+DHTTzKKn3tnty0pFIyhvzX7Kw6GpdUexqKkaqis
Sa1YgEl1HNF2jqWdjN8V1Scfukvm0oOvolYiJVn8/yMX8S6bHLrABN1wXmRKdj9j
Iv0c+L24XjggLm4EfB22nYSjaKh5WulVW85A8blozXUyOoydwWTNoyKNeusNj7fs
bVytGHocc+Kqz9xxOuZA4waJkeaxza8H3/gDjT7D7qNeFv/IcEcMYiqHmgQiIacg
OesKWZSzSC2zSuEGSk3CvMASJf5p3JgkR/NxbYs2hneuP5WVGjXDmBRO7c2aljZ4
KAmK56tN9TDcEikoSSspuNDCB/sOxUs/K/OxQhdphRgU72gYsewpBNn4Do3y0psk
GFP5fX9qK/ulsGdX5NmayGkF+6q/dYVoE+FDclEJUqplhsDQXi4xKtKuWthJB0Au
zmziRorA9BZhZkICwfJYcOJpEpQdlXicNoUMLBnw7bKzTGBQV6i+MMeUyQ+BDOom
DIU4K2nRAfSjly9aiRXRnL8hcvIX7GZ0GnJWbv7esGWw0BxCdpLBA3NF/1aQQT20
NyskyLya8gF7ZBWICXCs3yrnQoggypkUZqrlA+RN/cElQyxvcEWiVUmotlKMRGsL
rqf9PFS0WNrChFtbx4nF5XVu9tstaY21G4/NL1KrtaWa/cgvS7YFkVqBJitisZ2s
VlB31hAhvC28D1riZVSE3dL0t0gTl+qiO5MvDWEUSdJyfpuGfmu/4DOnJvR+UkQ6
bAcLVLj5Qrz+CsS9jgGJHhXBPNEum+YyFTmSJ+6wK8wNKz4MvsfzVCpQ1evetNDe
1cC3m9j69X/qPrFK1x7vLgDveCZkk242m0z/3hV8MSIwRuTwxoc6/smOaLqF3dQx
ONNBzpmIY//SH6ibysBkGvnY7fOTXHmxXqhS4YM0fCQF1FXnRmI7vVNgKa6ENUze
FL7Rlr7NEnzD4We+49gyHnZ8YSOJBXjK3BQMxiYXertOjlzNuvBriwfCmnuMuQTi
G8zuFrnk4P8KEsiRoeAAcZ/WqaTmEJXgQdircyJERql/U6oR5UdXQ8qkHGYbCOts
ySEeZ7FIOIVDOCZz2EkPmxCr5d7wYe0/YcfEYcXniExBjlOWmpHzUf6AbE3NK1Em
w0U5+iXdM1e/zyL7ymSaR6696iYf3d8Xr2rKxlDP5s5d7HZH26iScCABL7r0mbf4
L+xPyXCaCt0E2blrN8K+0gRM3UDyEB2ThYDOgrTburIP3I74snzSO/dIQZ8c/IAY
dqrTcvc4T0ETnF2ne/Yj2cCNHzTPisqOposR07Rym/sLG+547DeZsV5ceFf8XWci
pymxCZd6mVrZu6cigsH1iQc997UfLLAHyGmabzb4RI4W1Gfd1XfwcLpznXypxSbM
eByusQoTgR/3jB07xYxuyfn/L6JdYHX7HBY8OYQsvlWLeLat07CF5IQ/1vC/u8uy
9gLseHhF4RWlBn2Uoq85dnai7GQtuyWTL0rvgkwGbncZoz9+ZOJZ4UW6Z23pgijg
qZ++0BjXnoEtiHY4Wnx4kdfytMVQYGxaC8KOSmp680UmKVhoqkL31oDqysYPlhm4
I9bNPYUtlCSV3G0i+6g/KmAiLQrh47/ZM0QmgDxo1aOqqtszXv0Cj1rgAr9uwb7W
yZWjZyOfogxOuYq+wIHplfcMFV2M6ybxYrbDXTsh1ztRm7a0pG2yT/Qt/5SzCNM7
AajCQoJzuibiPD+kvMaNBGZZkNLLfSBw4WExt3PeO7mQS8P1m7nUgd3bJzq0DUSI
hBOR331gDTI4/ejPWXKyr4EMshnx64fmz4d1/YR6DAuSGJr+wc8RnOMU/Aw1CCXc
NDD1OXUKzUNaHT7TewbTZYhrInxZsHm6JAmXjQ/IoGOLScJwFon5PoFzviOvA2KQ
GyGBrRxN3MhkpyyKkM094nlD5mstVl3T5q0mFQsTx+tR+efRWT3F3GJ/moeLyseN
rFFY1qAc5YUKT59J3q1hY2neXyj4I4YX2G6DjOuukVF0SmTt5+fEyqJHkoGRfLmc
ljr13gt33avSsRLMjW/NTU3ABSGmyz/X5n8ZMvQ+LbByY0Q2n1X9myiaXyQ1ZWD8
Rq9YhU1K2NQeJ7hxfh3v6Fgdre+7Ub7ShgWZNftyqy5HjEGJmsv8muVATEidLO4r
MUAf4b0C1KtuukmZagAzCRtC57/to4Dkh0/at8gbx3mARbrmLCB0EMWSYB88AUOa
QV/pGpmkhprjcFzntbN90k7/b0renx9JxVCaIeZR1Dnhf8UzxsFq8ZBRw2K5lv1E
wCs0tfAmqb21qWKM0L87Ebx1tK85vzyDVZx2f236aeJbuX5nfGKgKeQEeizCNOLf
YVPZrSZtAs6xnO3TzJjYLktg6uoM8b4ar/KcfXeQk7on+RsZXh0154ACEZ8ovXw9
3XSds4UFjWa7w/LMgIMQ0fEyDIDvgSEzhWUEHQ8nSXAFLd20fAjv+/T7GhnG8ZNF
N9mjK+OsyMnA+OFvL3rkVomC/VjVcguB1+KlPrlwtbQNnsityZ0/72kGnDtt4t2D
XCtKMlqXFWqZ3jL8aavPA3SHIoyI2roiYxGWp2eVg0DxCtRz+M3tJhYXox+C2iTZ
5NN3ykas2d7RG1E2jVJJKvz2QlDVYeXQWMmMtkRSz85jSaz+4zlWltuIbFYAS/+z
brloH06HOuiRXErFLf3ZZ0TUAK+UYQsUOEIPXBLC86rgwF9HmY4q6SzW7OQHKfun
Ew9sz8OwJsPRkQz44aDVi7r4JGeVT9t7xPRzyyrFniMy4zj1khuotwwL8XH7IzmJ
/UgeJhUWW3Y2vI9crPtgrJ5AT8jwlAH6nPXTlDR/Uq7SXDqq2c0VW6lwlaQGCXnx
sPdP+rtVCC9aL4yNDj74J4cRVJKWhvksudMzm15yg48GMuyJ24su1ViEHaLL9u4b
TM9LI0Tw9o2cMdZAS6vowa7HsirxjwCxzM2niJwD7op8QrRbxFNyyhdi6Vj2VAMX
bzRRtB9x3+IyfI0NPU/vhBq1Minm69l+l1ltoS+EQbkB5S0iY9KtfZUN/BMY2r3r
uPOMdwZ3FyOOtyP5iKf+Hui6NSo8wrcMO67mu9W7tRkTtmsE95FS0zqkwAhYqGD2
iRiRxSvKQB8OA2GiLzJb6gy2FFHA2uyPkq5RaVGIB2Vcqi8y3V1qlm872Ah/s+3X
RIBeZGMTQ4yXB+zSUS9imBDKQGGv6II47/siMBEMZPIgIz/mQV+FLDXpYfQPe9w0
pNmkmPAbVutD/9xCVx/rMRtkqfegL3PF3lzR2V5VGVoIfy595OIQCYhVZQ0onIXu
7kllLqy+aO3sWDLnNJVWAZdflPoZ6RcWfUhmLEsUEg9taoNIQ0h6j+VUdZNbBcpp
fC7eNixIc+wRBQ7mPkVCUL5EsnOilVNgxBHOXzf3+Et6ZLPE03b9vZwKX61Edk9P
TJ6+mcmg1GicL77vqUXkoyo6yI6Rffl7AWPIILONH8E+Cj0w4eZgjL0NFaH8Xn56
6pBESr7j32Mxup1dLAYIZkvv6Vi8rGWa8NI3i1JaXoed5uhPCynV/sd6pmcndQfT
a6cQtuyW6x9ZYTdc0cxT/aIodyA682YSCtyhoQ9zhCsVmAOngTYQB0Z6tAcm5LE7
CB3rlNkLk8ZlXthg+0jV+avD3Y0u+SYBsXzr3uX1w8oDd/zMmhLovYWkt60/T1ah
NGr58B0wBgEeb+hWiPUDmIlTz5nLLTB8LVBq6nDxIlSLUN26TGRFyJMWgGHyDVqq
EVDRqHedRFaEqsMex2GJZ6NCbVRVqnnUg374h9+rtJYVsWIA8uhGQ5BUiNwkMW7T
WKJDFUm81izzR/BYnCIX8fdatMww8V1uGO+MTq74kgJFGQiVNKEGDTeelw7R6MAe
Zdmo0RXsL6huw3VDCJ0vp7ssoluCFMW6tXev9XDdNEqpkvRyzO2Sv/GqP2BjVWBm
v7WkzQbOiR+YTt+Io419L8mAD76qkTIm4qpXjLQP26SGXqGPNNXS20yuccwUZjUs
AJ2mXQigJfK5dfbtJDFZEWqpa0kNKuCUfoaKcx6R4dGnMW7rcdbYW8LuyaFY1zAG
s0McKu9XpPAOtO1btCfqsiGDLo/qM5Jp6cDLHzFk75bBIKbWUb2lr0NspmttL43X
2kxNl01N3snHEPtXy+tqBTuiJnYyf1S/HS9zZSr2HVvAXENKHt/3jkayug3ZnebP
RuyxdMmwNtcFhprVo7kwudwJO0rj5vEBtwLys9ncI4Hn7F1eSYviSHioPUfFlidv
EwfYJnA4u1Mrm1OiHHUFQqHHCgfdxlHf/uR+cS7ZZFsjsb89Iw8WkyRRj5s1y25q
JwoNWiGmMP06zNlfGpvUkKjRdynIDa/O/kIHFPcDu02NYuL5i8bDnd5wxZi/svM/
YFRRt2jyQFX6y8Y/0IW2JRAAa/dK9Fsea+xSa4lVoZqTEBT0bkugXJbt/GNE3tha
aJR9nVL+j1X3i9gJG9N1LbiQrPjiO24O3mondCaXzREOFAiOaVsAd7swaU8kZOcy
uYgGJ4N+/rxgYi14XG1sDHZXayA2vrsV0ykjEWuOTN0FLF3yydQSkBBR70xoZu2s
dS+k3UtokBMHtn8x0WTiZFJMTAbpEqRBSqJGIao8Ffzyk+Wg3PIgHR5gr8n25Yuf
BKiHGUW0b6+iUj/tQN4R49dcGP9/tBAM2YC95G+bQe7SONLT9lVfzrL7FtRfocKN
lUQ+QCiUtLHV8Dbg88DJdjeAEb6Dd/I0N7wddCFRULRp8AIPmfIhHIzQ8WCWEaT3
6r1/I4Xaz8bnzXanUOoAcWtWJT+FmBCY2Vy5UFlWqtsPRxShdjALX4Itu7t9rPri
2CXng39MQdypoqsQcr6LFpy3YUamgJplkQ4cvAjWd4PloOFtqndUPSVQ1/WNApG3
DxJ7YRGWVhAuDi4TWTGz4B9u3D9cLLQH+IhiYO4bbQ5W4CdOYL565AxDuBFM71uW
JxQuXH84jtKRHN6urLRdpGlw2gq9DM4+vf01a9Hn/wMrBOzyqaXc0MXx8SYAzw9M
zixOce0FpXsy3BQbzWuYgDgNDl3eagJohSG7iyJrAf775aGzUAKz2YdLoAa6U52C
Fs7MMakca+hPNC+y58FocbfR4NZEYqyqnACneBmO5rllbO/dSBYx+W4IUID+/Yls
Ai2/Lce1+p662gb9pB47Ng8/lTiX0fg+zOQC1qM+5FrSU9BVOdSbIwG1K2Pg8GqB
KCnwabyvnBMvCGqt6Tq98gxTC6zJvphGKW9jh0jck03AklEhvjsaZG0lCzL+n99l
f63b9RceABqSeOORfR+dB9Yn9UnHBZxxO4QTZBilcrbopGYQqG2+hUqtq8qfU434
OR9nE0lfrosOb4rBSQnu4n4QitA8WzpkvgpGkLQc2UnnKER1EQrXMSurjqWJ3ACx
/YCdXLPgrGRMb7XAlryWVjXJdl2u3bWGbAXR5AmkeTeBCjE42tUb6IbJfnZ0oF7s
DIpSfPP13iwHkmQ7Td+CArAPw9VKnA58bpRPbLcHPXfUO+xRc4dWiPlpUUABOfi0
gg4Zq6rmRXyDXPjfg8LmT0kcGQQZxPMqOloPm77kTb/EXpT8RVFrcNFSgsYWljlu
zVrDqHMFANqvxewUhgALAc2VMX6ljq4h2+1493XRtBA0iYKGFFxB+oqtufdIzHs4
EkBaurN8qxPCa6EWwBSy7LDjqjli+7jjxM4LUnaY6yD64gW87hU1mQGj5F0CEbvK
bD2n+cVrFhALn7gDqVPNqTLJLSdX1cfZ/mRgEmTS5YYCVzoJp+JrZeYhlCHO4NSl
hGsWh8uARhKzfEd77GY3jmPcVc8vsHksxbR5cL2ScoH60+G5G+xPoDxvu4RoNjQr
6LQ7zVMjB4k2wUCu81dQaOwDRuQn1iWdRvwbiKGuEyMru1vApL1WXzMrQ574WTuT
eSPYI5EMuDT0R0vL1eFy5ZqAoSTKj5SolbjFsI4TSeYRV71aaL1/30Jipq1zQ6/U
bPMFLjtFe1YqyPlNXCeh8h1RafprdWPXB2wsrX4LaduD25mZLsKK+PB6pC/OuYi8
vNoDNPFzp3s9g3EkJHy2jHuC76KO2WGQdjBRIh+HhqEvr7nvIXwf5L+5qYltR912
sbrnCl1NDLUIHXPnwkp7ut6h/A6wS7EQwWf+7FbPmiYP5xx8AtNo/oUvOVpnos2k
ffF/Qw+5jDYfASwZNQibYBd+Bgc/HTkvdrAEqGyA8n4AGC5TAZTN/9XZWdE7rXtl
5eszKutLpKX/ZkFqCupRWBYymMHUV4VKmF5XwuraHjF+qdB1WW1aYSrIhiRvLkkM
S+R+ue05gAZIRxER6+YyNI6+keqHS2n9Ls4a5wN6+6zBpWrlkXmZNI9BkzGNqjSE
NmuCGNd/TzfPMqKjbIZrWI3va10pyynBPElb2p7ewOBYXX0DXVzAW/6VRWI3k7Ej
ZVveqt2apotTm+YkDwM0nK0nCAjeLfV9DpmzPYRwjAcys7/fZUU2eYfFIvWV05mR
Vts/6kcreu1y04GDE0jTAoTGhGlA6peyqLNkWzL2LgsNfqh4WajBt2xLSl4RCP4w
cJ8AifJJVhpJaJpWauVi9IdXYAABbO5ceAimGNLaKfGOHGgtaYk7nUFtD89xVpJt
pkynvPeWtXnZt5bXHDUtoG9SHtBXQ0hHspzS6Lcnln3B9ydUBQNQRStsonFmODTH
yl0njXYs/WOWSHOGvW7NX+wgx1WZHUTKwwiVHveittalSBO1DcE+x+hutoys+HPY
zFIFchftXKq2NSfteINKr68CsMN0GHDKPUYj8fMgvWTrWTEDVW/K1lCiqfKvVEKf
r9RHrOA4sjj5P4F1mcDAvkJG93hZiQ8YMXOz+bl/9Sj6SJKvIO+g4hMKmqdmdLoR
GgkKx7jled2MORwJjpSb9vigM6i7PsyXRqYzgC6YjlZdaRgbN5Cwj+sa9DTL3vLB
Zf+7A1JFSV46BTNhnA+h9k3UYFInZloQe7jGBQJDGrhcctkDvFN6e+cKwrZsz2Z1
GW/u7rlMmqmFZpo5hI/NSv7HW2AQTexgcpzo+d7nIagHBZsMGVXl32nacy5XNrwZ
i9k5pYkwAgIQcD+ZjVMZRy+beO5NL3UsqnBIT+F/rvOxPvaQ+dkVUFnRqWwnynKc
yTJ+cdYSODQfIvLpwOMzvA3RcCHbRu+Rk0IaiRrKFSYzLphshtH/pa+PQIw8wBtd
4qm6TiTl8hGxMuUn3I325kNq01XFsb1n3AYG3iyf11znudGYO9U7ZzJKpIiLvGN1
QGyOUVsuCIFeSbaqcQV2Z9XEYdJ6GNQRR9smBniMcbrBs+QcsnHFxgG0fAboHgOs
AEeaq4Kx7+PH01F6d56FXPH9rMrFcYWBT8i/EW+7KjGyrAVTTZBQE54dLXkp8H/b
KFSNfqFrnJAkpsyLFrTEqMQivjbwFDmNgQfTyVVcN4LzjAN6gvoXeI8Xsi1mrJjq
ZJkYccjDBEDx4hPY8SsGD+tzXdnQ33ItenL2U8FJK1exXVPzAvtIqJ+FrUdTJJUt
UdN4jF/aSeMl8wX7+0LuwWw/4hBF8+EFoE+u9c7DTP49ZKaJGzu9TQQ4jmeLQiJ5
bBLw/yKiMm/Kp627KGr/smmdqnynocXR+FHH1Mw+EUy1IRo8aQdnQZp2RcZLhMoZ
rW/FCB8k88EnLbFdHarQZ4Y+EOAaR6VE+/0crq+1HrNMoet9xFEq9uZOrvktxCr+
cPd4hXT+24Uj4tQ4gQybNOunsPX2ZomCH/uapxWbLK8rzAut1m8eVs08uRUuR6m/
ttl+OlzGq0GPQyGpbPciiExRYtcILYnjCV88AxnUrsS9F6a31R1rENYk+rf2eq7x
DUnmFX4T2z2xySDxbi6EUplIEDMHMCYsUaQ1U1eSYoFbKxgpqsLhud52jamelYWd
XaZRjgNuvuVi1eCX5326uxOWZK+rlmD0VfqMnplTAb2dBpFtRAdzj2prSRh8dfIC
0tllG+deumAXq35e70VSspWpxAYj9Fc9wMV9h8FzaasqKOr1ioBIULRFpIPgmmm9
kCyRgQ0G8Pbz2i2FlU9RGRhChmyaEbv7YJRlB23TZS4E00uog7SUMvVQ3EI6YhqL
adkvf0ZyeWBRgW1YQmENaJCwiQNg52ZNS0IkOhjHsDvOyijL74UvZcaTm1/jbV/7
CGSChu6qaX4QJbRPlpv22vF1630tw1fJuQ8wI53HeitUZIvq3ix5PaSaTFL5qmxM
EGoaGTZomjannO6JMOQEokfHIQfLHmGvCjXtQSCaYcIZlh/EFhmiGr9XdgPWmT0Q
VugpSU+bLWFVId0HYHxogRJhJsLUqzhUhDP8zDK/api9pzEd0RUEMyg+tvUYsYsH
BlWXOATHwxvJ45wwpG6TBEdiWTrvr0ozMBCOLxg29JVssPES0Y4xUzlAP1XLk20/
vapioRlRFKBuYsLpE0Sy6CEKb4cBJpL+ZGu9stGtWYAuj0UK3I9c0QrmAWhoXRK1
8KyWM1BXPn5FZbNga8IPb1c8OPy09peguXvXxZEUPPRIb/nn2QBleM64xj40vzUv
LR8KbnBofkYho5hz707kq484p3zKHaVZ6CpKkjNb+IQCc1/kF9SZo4xkmWguFZ1z
PsIgdoSIuIma+k3p3CMGy2rmp9tsJHweo6Y0saozoW8AEcNPDf/2URWtrec2ndtK
6Px4EGgsCl777AJx8yEsWGGTUOYMr8YNAazZKngERuDX9CGnoEcPyQq1wofItGxN
B14QAZwi+HblDCC8PfeEKKySNZJXeJhIMGCsFM4pbjVKd49oeGoq1jfICqBs2qb/
hD5C4Os/cE0SNk5VKRlHQ6Ub3qy92RXPe4SyYP97He0/8QbsML0yhwLjTMqXfSre
gFUVvAVq9qndaL5OAihxnoGhLrbCNGTXqMEyaFiLN6W4zWv1PZL/JSRUpQtPxjt7
v++8yzIbi34LXxLHPpuEaF7SLkvTMBJEhn3kddqWZbdxANMfhw3Xn6vlMlkvTfuW
hI+H9PJ8eZcSSYdrlcNb81yLzZ0jlFgbIa6/88vDsq0JfEv45uhjzdKA4FPoxd52
jVaGUdi2tisZT2Ub/IQKpFXJO2drTKUI2kCG4cYrpDVkDyGHG29yS2+mMel96hOa
azIQGPJsCsjjkD6oZEiIRpS/OETkV6Wl8W/B7OQJodNoR+RR/J005cuVZ8cjw51N
whHC9g0zt1/G2I+yFJwv97zc4VA7KHnbT8fDKRuMfKxuostL6wUjwHfS6yqkyT++
VPoNqJxg59ZHv1qJS9HtrEVwlEqKfUI/1AkRCd0xpe5yd+jBv6tIiWJ2Mkpddoxk
tKuCaIgJdUb8W2ghTqjlrGFrUB0nDChdexl/GZeB7UcJbBE7Ew6JipX8Lvx5cbBz
3CsPAJ9F13mBApUScZP0ikWlcJPluYJhQsU40ZNXj3jeXjFZWfo4TCm6SBtcXjSV
cVRj++EUL0AT2Cavl2hFI37kF1GwnrMg4rXPgmXcdgnt6hIXjadlst8nI/8IB1VN
LakfeZeTNlCgtPSmngV2Odxsp1ax5zE0B+VNQhBxITevV81JW9t4C27w5e6uaQlb
GMxdVSo/gehdPoVBfxUpIgl8htOrNWV+eA/9hLOvGjiZ7jKiXGS6FRa92lUnv1rm
VkGVr2fVVEMyOefkw89jmawYqs1UXvVyrXKYLPAUmLXVjm3B0wlzDpYd0/9agfxP
03c/tvmsludYMN+p2n8XkpF6RFJs7Pl+iqzGT3QRROmGz7L3Iru8aygcKfa7LRtQ
11j14JMM9KVtQVVAnV4Ecj/GecL0BlLTpeDO0LUJ/OvFVm+TURYyYVJ2NbFa98ff
fhr1WzMmfsNXn4lHlMdvBhZIUHZaJboFfvY8Rwo+BOkauMg7MVNm5gCiPN1sjF36
g8vYFxHQn818uk61u+WJfv6bmOIxHRu4E+YMxqhI7nYFrBfF3qPZCJfrOI6BVIE9
P02Jjj/+3dte9bfiKt/Nbkzrn/6lskIQEPIxWZhcMT/gNkArJ7yE1nw/Bz/erF0K
Gvn+4oMVrQMBp4vdnG2UwHEuoh858r9rBFDh3gjw3eNiRBz7Dp5CM9ztzOjcuEMb
DjrdNVBQxutCq0B+cslPUHTfwIVHyp/u6n5T2bxMpxz7MFhQpDVvjiX8t1h9YxdB
SDl9wyS3vUxtV2rWIGOp17fo9XwwVo0AQLqZU/T5HAu4jwqqUJ3GD0xzZ0hiQ5Fl
Bmn7mYnbpG1fVyziNM5SuwvSbITwBgcg8739AqqHoO07pG0Ua2KRLN60hDoWl8Bx
ATBfflzVYa5eP2HQBvVCtTGaLQadKorTxgr0jRtXNSbMMEE6cQvkRHvyBkqlST93
JpCnNEklXeLCNwTKT9qL3oy0Np9jo7xoYD1XL2AjEej7mKP/DStdqRDm1RWJwOhk
HMI/6SC9+UrTkTTBDUgDH1zwbiNdm8UQnGv7QxpT1EQFY9W27HeA16zN3wvvS3Hl
jbqOOIow/cXbTRq/Z7MZ6kt0bZBN8eF+jpFBUE5Fg9ebybpzbtWP2aotAZXnCkSQ
eLR85hioveqycq3Lz+Zu40/NisbordqP6xIgO44af74tNTPanRgNGYGfKcdlFEGo
+c9XwkjmZRIzpCQngemECG/1tAfs9LDj2IZ8ISUQv+hhKKgsIjPODX0q68kCMhb0
PR+lr32k88eZiuf/j8K3EI9hxidnT9/RDqKOMdJGumxQE6qmb+18bXx+9WISLqhY
GfF0SrUC0ox3avVV/Yz00e3qDGJX8ZQgTKY+tG7lF00CQ7iHeSFqIyyScXCmr6gm
RLgu02aAVHHgR7pcZNSEK+3gYZdkEu1X15wQsqQw0HBZc6w0a59xxd5Q9b3W+lcE
nkh8duSg0cBdQCuNdM2SF6UXjYPBKe0SKDra3D6NJspayraPv70j8zrSWURQo7Hy
LqZlkqc4nbC4aTR1uCRgNBJKFCLxCYvC22W2CqSDiGyVtDnMncDCVsq/QcqHGtaS
fj5I3Nm5sgMgMmDLJm6Il1f0zpbJ+QICjxd9L9q8eZ/H31hw/grJ6m4tkFsmEiEC
K71flCup6+9065Hz5+QXdVaCi/prQ+i4oagmOy9TyiJ63B6pnVVrLtwDAj8I10TN
jQIivn2p4tbuGl95Em5VAitA9s8h4nzUi57ucryJ4Bev3Zc/lq61nLYrpRgkqOx0
PYvtJt8heCD81yi4F/y8cS+araMCA7bHCwXX+sFeS6xKg/RC3EJdR3nqOE14DRZt
PSDjzC4rvBHjgH+LSCrLtYKfGxKnQd4lwCy9UfqsMt9+eI4tymkWaaFmK4ZcZXrm
sytAr/dIyOt93obEpvUsDm2gI3s5pRqXmzdq6dl0xr1121aCHQwiGqD3EbFhzxCE
+qJfgoIGIOALLrROCFVioa1Z0APrb7vlezVUHH8FuPdU3ofz49EISl9XqrKCWs2e
M4mhqYgnrT1ZqbRsBREDI8LM2AgyGKvYlS1noyc95x3qVSmTeIUO3eN9Jjs+iZ/w
GxbNDrWObnC3re6iLWFjXwUcjySOK7ziBnQyEAPTlSTlHJpZID1ohNErtW/89XLQ
zQsWLFok1r980glD/Zo1ZaybHbwYqic7x61WifLIzECpE0uranOwx7mOVGr7L31m
E/jJ3J359l4NGhnVkLMeACy0DM5xptyJK7EFMsi4V9Q5iKVNSXJ/TbIJ+XBYVN+H
JENJGcLypWLVdgoOad6ZYAQ1k4l7DDi+kX+Lul2jAUtSJNQmQM52DlL41581Ar66
LceoHQfC0Zb0MOOPEG7Bu3dQi6Ev7sYzQs6O8JBy3N3f3ZxNnh3Dc+cgMLM2Puvl
O0TfJvnFvswOc200yraXmRwmifdqiyZivgM9+GmYaNGyOXYGpDX+hObgikaml8X3
b5achOl+Zt9ey0wLCC2ey2EYolJQxvwGZKi0hkbquXLuq24SM0UXe/ZoVRMg80Tt
iPLRHI3/ixQTIZRo7jBlJoDUpuwvb+8MNHkXflWo9+QOkoI5SKvLXN4jat0Ienbu
3CFz4WwdcIeVyXro7b4r/2JILK6KoqbYYdXaWNTkAivIJJ0NMn+pVhnVsMGqstLh
eAk2HsFi+MBc4t/M2zc9jXRVDrJzOdH0FMjXkS9s1LyO5ephCVBs4oI2YGGkwCbW
rYsVKwnuvXrKP2rniubVRFueMSlF8klyAHdWGpux2w/UcMs/HzeEQ/wOWtbYetCB
d0Q050JIMKQp3WjzIrMNxVIbMk+7DtqJXqCi+kmRHKxe+LNPsyMd3jReM1LjGbQV
QD/afUqQTd4oHTR1pa4kpuXnAqhCNjU2tSzhePlUGm5v1f4DvLqCMFzUOtAdBTUg
CSHfXtgRnH603yO31KJCa3louBdmztQR39lBbycTSV6WU9kRe28rNiUSo5t33cFJ
d8xojaGE6LEvR2u7PYisoiGBTiaOpv/URVV7dMGlc+dr7yr44HX4LbO/mQR8tdRR
8dv87ZS/+Fb9XlAJYifJnrfQrxjYIH32K4u8ajS2Dd+QdfT2eM057S9O58DLpF69
CxqA20f/qg8xhSXBWAW+I3OdGT+Q1WIJQB+vqXCl6O17zR5fKxGTeFqxOcQ3LazX
NoIfiXBZomdqBswxCfeRW8VIDZmA6syd2GxztE2p1gcqmf9FAzP83PeBCEY4ogLB
+CEqnwMN14fYqYRJ9BB5ZCc68uVWa90E7Jq2k+Ylo2N9RzqSS7ULbJhOOVItZSC6
f6zlivyl5PXnKQCzA6AttWSCqukfQIX7uBHGroZhtRalyPPIptFCQE6ViW5V+3/c
g6YTOLRBUtxYeO56TcBYzlFWnKEtCRgNfqvdw2cpGtbDMCuYwthKbVzf7RYR/g9q
NPfdw2vzi6WBQxZ3H2vC6qGsAi64FxpGoMPdMzDE9RPHMSsFughUpXVUBtdB3Kuf
R/wXW1mp7YleRWSiXPZPjri+rufIKiiIU0PDPOhMAFN400vmvElqsX84X5ZmJTOa
hmqFo8uN95kX0tjcvNVRdeyQ+96oCHfKvd5wS53LYjbMXpvlcqpVIm9YLUR6GwqN
OkG6nvYBpaRHqCudR53u9rxTY8k1vF8A7a5gjCjaaB+hHs1f9Nsmk1x/M8lEf3D2
2D9Nq1ZHgrYdIcXSbOcCvjz+eaMBSgoJ7T6KQEaoC6sDLRg0XiEQQ614JVOW3fh0
033UzuWkml6UZkBoB/pkvQa0h03c2it4vxb1jRXcci8U4rzn1uQR9doCnWdWz1y+
Hgh1jrsm5XAckpYcJKYrYz3tKeyAA4I0cOQkUeyXkHBibw2JLHCHMNhHHN1iHsfb
/G30Pv7r2QX/cmaUKnLBOUlnaC5wze4YSQjmBpTF9SqIzsr4+NwzVaCltsQC2rTD
BhdWG2mteT0SphyKGHkLndBLS7g5QLEIsyuJAlHH793zXTNfAccgvC7exZiH39fK
r4YOufCA2Rki8Reu0VaSArz5HI2AqKsUlf0r3LtrYzJ7yq64oGxhbcc52Vnc9rrE
2X1NDUAmRqRqKR+z9yKl5Xas6/aE68hpp2v5bVS09L/pzolPA0odu1OEXml+oKbN
1WKRYOeA9QNb/u+8HVUoTd0pXCGyGabDRLD482eZsuRmw97XfD+0wDzEXUQwdMEZ
Vrobzi5dxrr6G4BKm8NVuXZSbFUZhOnUvkkzK931O8Zj/9BHDT4I17RMktCllQSZ
9e4A8Ah7JFX44M/lIQvzMIsNfsXm+ighC5m1vvSO90AIBBjbTZ/IIeJqzh1ZZDBF
U8ZUv1s/+RRiIKmlGv7MYT7tcVxPAJYDcwSgYxy0AqI2oWDIQ+4OfhtD97ear7Bc
fr7+29eyaPyU0iWh3Ji5wF/cIhIiDZ8nA19pi89OpE/xxPb1db0vk83Rn4uStJEz
9PKwB0e7LvmN/XxUHHZVj2XHDrABz85jXPES5GDRek6TGxcMqeHTef+f6JWY9fQk
AMh/fWBvMSKAjNJ8KbcpLl+HgD/ap2UYPuYp4sQMVmif7t+WSz75J2+gTJkUmA43
xeEBAplzSiBL4AoVTsssh87tTvBDEtnRSW8/XHBa4i4aiPATzc7YaxYPP9lXsDEb
MTXnfJ6m9hLG5THudmL22j8Qx08BniQT4YedHTfHdWK3OYzr+P66pJRKYjbidMBJ
jNrcTvg/mB0OrWh1ROmb06XJUl6FFxx5mo2A3JhuyVaigT73Q/EUTsMl13Cs5CXC
kBzLUa2Xsd8SXGRVb4jkz+I2Ifi2f6ZKId1bJugIYA9VzqRDIwsuCoet8TF6vW6j
su64BpBFvqkGtOa7w9LVskBBAS0QwMe7dcdsrETXhGiqwGVQRxPWTNZvgLaVNypf
2HIY4zkEl6AsPRTDoM6l1o9NDGgC5ogi7hVU2wE2MpelimmGJClIFwNcA3VFL3Qu
MgmzTPp0GuM5JhpmoC/N1jmYGeaCvH7EZ8W/98iMeBehO+sigU2J18RBUVQ04fpz
HqimRIzyEwHmJYjpyvXdgD0lU0RuxSJu22Lh4f+ejena0STzWiZxal+FHKQhTRmD
H3r5bID8CKQ5i+bsih4gP1/qLtYapA/Rg1gRru4fV6p6amY4Z+DgkD/q8JiOIoVx
tsMMfZA4FID0x/D6WLUzsv/5pgJE3Qk5jSC2D6/iBS5P9l+eSt5+iZstEsuEZZdG
EQlzIs7Wb6Jqr+F16tsvFMAmkz7CCleJt9r5PEDttH58ZY1eZyatnXOdT/k0Ta/7
QzWzl/8beSJzUs9BdmrRlKzSQM4TGvWnha1NYv73JF51gWmMph4SYMcRdd46vjP4
ml1CkKjZUMgi2/gYTIK9wLLyfoPCXTcVVxhNxVHu/eYGl+wLJLaaIMOBBRPMnMxa
1VrTxSjzmyRjbBEn2jc0RLBrX+5qgbmpWI503K8sgkpJo821F/UTZOSIoZ6Gu1lW
pgsffWiWxIXIHfz1ZZuGeKMIJ8/WoeqRgHGjZWuHuOjWa3S6ON3AIMEdR0yD/hKK
MJZT7wZxHeeCFWLkGC0YI3H7yaT2zPs9bXSUctEhi/lMd3f+S2FfyrtxQPh12D9e
NDDGUwzS0wzEV1yQIZGJFyI3rZXycyjMngohLPK3dDYaeGl9f8nyQlDX1gZyRf2U
5KI//xvGnn+1kpl7YJhSC+MJxC8UsOPo4tR9U+S3v/q+bJNSO6GE39rpjOUKBsuu
rQfTP+NTBteTse4Z/I/ckAXo5YEcb8AFoDvxSJwxAtuA9W7FRiaQrArRUtAOUZGM
2OJzpeMhZi71puCIK9TMXYBbEMz5BnSuDfwHUOMM7qCGHTCN7qTuZPdp/qMyVEu7
bJ+SPbbe1kD1TCP+njXz1kaS1p0fv15BnV2q16KCpUdJnU3d86sxsnMkUgPC0M7v
vbkYUcZ6MMPgE0whZJKtfZSDrdvwpHFrVsc1gscyHbvChqDNbMhC2OTSCjsxI5zF
VjpfbuQ0ieEl0/9thU9QSghx7CAj+8REVoq7fwCe3ah0S4tIefzxynEiM0SdNxZK
tJ7a27008HMnzC9FegY1PuW2+90Gdir/kxToNcARHQquy67TKomj65ZWOVmavEUw
oVJul8redGGb8fFq8ji/kkQHdTlkrHDT9WXtQf0PWRCKnnNBsSsXwYILy0vu8isw
HYVTHCp/qc8TDnQDPl0qvQLJ+yMMVR+bYqZePBim+g4WOI/Kf1Y5bRZaCTZicOXX
F0Bpl1ypVLk7v88zlB0aMy+6va7UvKroa7vG1/+56WrKE9N+NttktMqiZIY7J3mM
irpytOPDRtJ7O6X8R/VpIAyj0CAxHtKFFDCrhVcuHhPNyMdMZbpwYhRyc4xlS4RV
Q1sCMYyeiRNCqmx8jnTKVza0nx7B0OT3DEnf94wLI04Dzvdtl0uylMgI38OEmahP
zyWcUkAM4xqBQc5JkLow/iiPO4Ay6qFUnRmIVSX96iHjoZLcES3ZNw+I3TobkPn8
QcuxSJq+Ubc8ivF7azeTSZ0A3eevFv4wqPR6WhkH7LLasGtvVO0ejfEjJWUKV3i+
/4qlGLSGKWOvoio2I1W8dI9tJvM4RCdUmYRVEAzOWukLYZFUqQLoqPBerZXSY8pG
TXeEwpqpj/Y/vXn/Q6qITX0fpYOuxKtFcSFnNQ8wXvKinE3kxwI/xDqm7vaeYBUP
cSp87qYvxLr3znGzH0zovEWpkE5dNObNRP20ZDY/zMyAtk/rMehFc4IqofHS38DT
8gRfZvRKsHzCb0ipVWpQnY0xWYk+CCLaigeWo1eEsbGLCB1F985vHc45sGn373Gz
Ad9AeS2HWybtFFadnvPVeGn1lEDFDIUxZ79y3HHUYW9lsdruZiYJ2PrCfsxLajpN
ykOoo5w7Vxur59q5xfltEjPMrGZlW2clEobCfss847r4fOMDwqXs6MTP9IR33aUy
ov9HwjTY2w3USKFXUNcS+msM1jI8I9FVjML80EKTRqaem5g0mRL/Y4BjwCtNiCKr
AiFp3FFCXHEa/mU59/qyq4cu6Wqwt+3BEvBYtLORrY3bgseJwFBDZBu0z1/p/ZWL
4juSoM1X2uVwutcFQMINi5iqGenDWHfyrZjGUw9my2VcGYTDNKYL/Vt8jkygoQr8
bjZw2/vvKrfbVE4FIPSjkJb4M9q0ZmwwnJVCrEuVFzJwkG7jaU17K2jF8hxiPb4y
OVJHpodDooMuNWzpv60v1fTCDdVcaPZveptNG1wOC2XD8zIE0SC7xqPzSZ05GFy+
mMan+Pex8y0rFgfKf3sjoKnto0oufvNx9dpxK5INA3diN/OLIAxoyNMq0eGR/EGB
fGLQ1Gr0f6Hc1/zUHXGZRjpx39Z1tHUCn5s9+Y2fer+2GFiPbG/m5eVlhI6DUOpe
ZPpMEpOGpZZ3vPyBppT4nCsFhfdzmAaQ2dzgGZfAfNacyhF47bzuOQ3YWMvjCOhI
yKmNc6DiTfadlWGozfwLbMsdeRTshXhO07QOlpUJ0+dwuJYpY5Gzh2gFFbVLbAm0
O9EMEU9OP6y/F7ZCA5RxkhqCvY9PyLLN3RBUa3Lvd32kZ/pxAeZELFIx8PDgAIHx
ul4HpL2VOoTegELn9BdPayU1CXv8sJgDi/hihy2nAH6WbhRqYP4/XQTN57oT+ynH
6Y0i6OKz5bZtyCmIoJbXPk2SFOeVYO2zR0orPWM1YhjiaUpkebcgiKgqBIkAseJq
zsRuA/P0Sq6bU9I5WzkaJTtGBP5/6eVmRYEPjqQSlc8eBO+y9btgriaLaIMMS36C
BLdHAE6ZX9oFFWDgZWYW31Fg8nDCfo8paT4vb+NdF7jNfOceOB8pYA4hM1oxRFwh
HiRPC83TLth8yfFvTV1GgIudeVC6jZrG+01Ns71Q87qNzilHdsiYSbsepwpZge82
6i8KmILmJP0LeN4eyP0Tx+1gIQar/cGbBvaH0eOtI3oYCmqReOT9WfsLIg0hQx58
Uz6FVmPSUlfSWPvKoq1H0ar96retYaWE2MLFnf15Ol0tUjPNJZKS+ll1i5wwY2vP
wNDdux/cHVEe1kHFJ2fOA81w4uYrkYBZWkvnXz8iT2XbVevWlVFGlSv/OPgtMi2M
sqDNnt0gLtFzRUv/4LybbDQ5qTJ53IEhCkNmgoR0mRs9QQNB3FycKdyzpqwzoh3y
Fhma8BdXJ3m4fei7KXGEN8wXOfjJQQRBYD0ZY1mKTOIAUY0nsjXoFZk+T1gP9FAz
K1Cc3errn99C7Znp1gGOyKdrWNQMg425ixZmnJeuXiuiYszJP//8LqnQCE5PglXT
KJ/mZ5jPdLQTZgm16chsf7sIZVhHFAH3AO/ApmjLwvVK751PmfW99DXfs6g+8fhs
PsR8BFgvhAuO2VMN7v+rnQSnXXSRAjDrQAzFKcAu9lzk105xsZfPNgCyfIK6GWxO
T4EEfzGVElAwCytmYNLVS/Jv5GQhalU5pVaeJD5NMJ2T/8PyowKzdQhNBL2/5KO8
ZIj+HR8ZzMydUlbymflF/bsJ+86AR6ajwTsDjJOybAWi2YI8z2fNM4tiY6eO42JW
disqxzxy6Cuaa+UrF6V5bco5itTcpufdATg1bH7Gj4FIHnfXcouNlAbxb8+yHXiD
T1N3YOhKPWwnOX6xjvYiAaMY6/ttHIs/jwKOTLr329ISHQk6mL3P+O4bY5UuJg7w
efCdPOJ1JojH6fjMkcLoK3ovRiMlVp3i1ILs/mQDiqGVyXRsTbjcmbiuFeK08POu
lxwA5QfEkf2l6ZYZ66r/tOwLcCYIByZdhSEbq8BR80JqGnL7NpMHvR7jtLDkn7qe
8bTLFYwIil0POIx6P+fQU4JwcUY1NcaV9GaRkT1+/+6xqIwvXmCjR3drAhsehuV/
fCN0vJtJJyriBXXMc1QhVSVWKAvt5Z7lm8ulgc2LhyfkFwdccYa1+34FRYrY0PvJ
VMrbl1cYlnjlRsmggt98U9VLYxuRodiacw0ea0O0x1M8sXBh89agTTPt2J7oHjL7
+8smgQ8L2ZfdbBnv6fs7t+LqwOOnvGDYZgmpJoVEghiVQ2sIQwUVAbXGaPAiw+1n
5vUU960CLI3IyzaN3G6MITKZroKrMugrlq4Wy002p6PePLwH6WsEHUP5k/Vrf4or
7L8WZX72GXa2XvB/rxoVWLNeAC8f53xhLaG6FSDafBRS9XSbxsim5dUpRKOrvQin
YZB4M0b7mli1MIaee9IOll2y6jXfwEumMa0jggSCssu0kNbcDfZEOTpeBpoHmKIz
5X1NDWoCq8z8cvEie11tanv1isvPIcBn3WyWDWXb+DVQYPkVfkk8CZQx1gq1sHPW
qKiG3Se70SkmiwiRh+x638AQfTtjVQIFpYBd0wm6/amriDlglj4kDhPPU+D+rAOV
HnUGgEgUgByjWoHMh2cr+xl+36bfAKPpx4+9gIijMtIzgNq55EIqbQsWFzYnQuvw
BnI62ZpRcS+NC2WEHWvJbXIdB4At2wyh8EEuXGPOCfRDYUJ9O9yZz/Z9XdzSvKQR
Od51BdJW8psZdRmFYwPv8CJmIjKghBk13pxgDKzav0oLN1xKMLySeziXYxpEuDE2
+9WgH641mMQ0RWRJq3Jr/zTJ6rm/ajT6USYdvSwmhK4MwWGATeBG8JcvLg8FQsqg
1dhUjtSXQo5yN4MGrXtu0LdPPd/bEzJP5rq/duSmEasloXzEphhXEusDKDHs41OL
TG7rMttJCw3+IPNnK2Wn2fZDV6righX0AU3FKH15fALcX3gWc0eQcK3NrbLz5PG6
eYrdPFPrenSdTAAZjPPeOqCL90NdyJe3KNdaiQYahpBsSYar1uxrv01CcAT5bwHg
87GG5h7v+d+YpZ4vMyEZbzkDza+5Y1MettetPtHz22YMjsWZSyC0l4+YIcIFe310
NzUBeB02vTMzht2YloKuhdHwvpQ3RFpp1xGIksrW0jtZxWaLQmIru3wibg9n+yaS
ef0qPDGBJ9epndCi+GeWmOn17+PFBCkyy4/4GhPVh3Deu1MVJevn82V0j4t4jr85
+qWhHtbJ3El9v2S0FIxX0QUGdlFDK06xxgy+3yF+YZrdijhXUTYjJhnjX9uYsv/w
9AABHAS29GwyLOQKVRwpBHBSbhg34eWJyJy/V045af30mFbothZcebGBI/0Uq5dx
wKDqhWpkjo54swlq5cvcsi3Bq+A/l91/gpeihng9yw9GH3nqImt909E1r2TGK8c4
oe1GSWpXzMYJoXE2yqyQMMcso7fqE1cAvYuJOYpJYCNTCIvMNVnwC+8IEc4HX7sM
4GnAiHE1B0OH6IE/PYHAUsFGxjab399Uyp5h8IHSeJaDmEa6DQr0UYnKbCv2RbPm
aWAs1uOzpSu6h1e5Ma6Q6ubqcLQ1Jrvu99cjmHQfF+gt5aGtR90PBOqAP9vC+gWF
QL/rJ+AQjxJxyjtpS4rIP/gDDGTQ6VYXixOk1x8kYQavD7W7i/9OLDtZ+Tia4/oO
+La5fNfVKQCOdFb6sX78XG0YjbRlKjcHZXeEWYsaripC/6/THQgBoSsTI7r9Cny9
6/VImt0WqTBxCKp4A7Cc/Wmfdl6PLhZ+dwVBgblEuqUHxeNTA1cYUxO/6slpjq7c
w8ONE1mx1X5mKgPXYbhfFuH1ev6eZLgvpEF3nxI37uRF/9pyfDDTkFdbyeQ0o1h4
vAMWrm4cixQmA7rZIIgbbI3r++dRp7yuE5C/g/2SxnaoNyol2+rhnAP3Uvpwtqkc
55VTlCJqSa7aaQ8YNFq5RIRGryZpvKzQJiUP1V90EsjgZQY/1ogE/dAxjnKt3eks
VVmulUBP0Fl5qyM3QfXdFpmG0dK3m8mHc7GevDlHvQcZXPj+z2sYVbh1CefKuW0d
WTzOG0J/myBdZeVxX5V1uJoIVsT4B5Xo2/7eHzU9Xs4uJIgK/6aJcWYmyxlh8ATi
WIHwTOLY0OTkdKQy328ecpnaePIUviTJ3ArcrtTRld4gtItdGCLur3kqtCJF75tJ
aAmviw75hsLpjoBO47JvG3GQW2ZZ+p565jdxodpF19DVKrq6jRhZL2LsesMloDSg
XcXq8/OqV/K0J9Esm3h/auuNhTIvKfJr0+2NAGSmk/XsXzd5XgazOkrElT1aFDUm
6NVt28Vr/yUKOtZsocd4CRylZV1Vx1P9vw/P6rLrEESVYp4Wq8cE0pIAWoMpq0KD
PHby89JQ+muCAmWF5Zdzb/9iUY/nIWLG3OX+LJ9wDZgZceVnokKlhPxw3cXA7Imp
He231UhE+bkfx+rs7JwzJ5FnG2yeHBQIN2uoEZ0UXkZtVpK9KqLnUXfihwiiRmIh
h5hvALXOkkaXPLwOsWyXGEiHSwvfi6ZDFocZisffXGuT8fwg4Y2hGmLP7PKOftMc
qPhXeHj/tlIy/tLpyj7sXkwD9A3aH+L9B2EqiThfyGIRoCLPknaEGqYUtt743o8g
/h/cYaScV2/XI3qonViPZEXEQu9Xsz/e2QGR5lFXFGmn/SPHwJb63eq0pnxOhl+u
oDTW0vcl2vAzWVGHHK3+e+dR2rj/zzD6Y9rmUuR8zU7AqzC4IESFx1oCgiWpKKJY
1viBGkXTL00szSb/Ay19AeWcqIQ8KJOkyEv3TVzVI5cuAq64ChKzzE4N0W+e2xdb
laaoZWySOLmNGPqvb4PbChUaL2GBpJr8GByCHRTntMdVTGlL4vWQioc8FOg4sBY/
gZfJmN+v5vtLzjLbqblOV453Nvt68ODFIE92h9AdPVcOHmoPjRHHAc/bxchnx71C
uEO8UTsENnYnV8IZCJMHLEM+aDJYm/9j0l8AmLcWAukxSkGiDgy84KfFc0+e//Ki
tY469sC+8dqFm5PCZfwjqsoqWbV+h3+w1oqp+Jpk/FJjuFJEWTRqewmMZ5x0yJNX
VaFgttrbdHd8mxiXwdY1Jqy+Nj8kEbpP5zl/Kksi0NoKQy8vo9S3swHMZ70flsyX
dHTPGg6ulOwot465lwSNInTmBoP1YgP432l6DBAQUEptBz3nq/DRKxS/akrAJ6Cy
Mu1OMpgDEqyQD6mYBFMgCbscBmQvxYauMMfmsnSxGxPj1C+5Ad0O/GswpmDbi5rd
tDjFZp66iM9V/vlbVcv6a4pzffFIVac0rZ3iC/enGvmspP5jf1bgZthfpDVVSA2I
8G4smwcID1MdrLjpmlZmtB7qU2lkRzcU4ROAzQD075IhZfTs/GBRispVaAlt16Ja
XK5ZzxWXNwvDWLL/+BA2NEseyXEudIK2scXBrrYp8k+mPXcUkgEUmSGA+MZlnrNV
C+xmRo9D4qxgX1/pyVBy8oPuAFUMhZ5CKaN/MAi2BbVkH3NKiWon7JDTx/xMPmdo
h5u4Hsh1j3HMkpQWQassiW7Sxycz3KGY3YRkc/Kmzthq6ADbSh0nvHviIAMFtjUa
yKf/0PCfW+erDiTFYJkU5uPi7hJ0JhpN1A7ZBBT+upkxzMsRMRJ6MXVWGypTbFnz
w88nWyb9K4XvIU7noNNivg6HYCpd9/DgQQfSRe3ENa/+HKx2GIn3/0aSHP4ci5zC
YCtlVZkjQcmUXxDBDi084HNnG2Is6McQtUhtnmMzOORKQ6K7zETAfbFT6DdwUZWN
y1uv5nF/4XNfJ80rZHCg6PWFvX26wA4fUA+hDEpS+CwPNkQAtfxuMhuZg6335QYc
LV+MhTdym9l7r4oESohEKEsl3lq69VDUD5liJAfn6ZalC0z1b7hcVTVnX0ZmuJhm
ml5fR9VFjgpINLBCKGVG7lW3BnCUf4i16QBMppmsWzpWZ8E6igj8fKud7ug8bR9I
xPVrKpM9SJMFVFGZ8uIM7nSHBth9iIOaMlot43NzCbA7cNHaSVXqZ5YlIinIlY5g
0xucNZCoC9kXACFd3kU7MNNy3X98lhQZXJ84GxjTAonAFmTI0Bf43SP5GjDenx2u
0WXv03L/wiDIkmeKSwAGIB85HNQRcYjWigHYuQhzz9kWjtV4ViecZBqqWTnDnyrS
ruJXAZ2IwkTy3NeVEOTrWf7kkpufkkSVxJwc7Ojxt646QP0T4K8i7tt4OrWlw+Rg
8nPtC1BYzp7wdtmR9eLXF5ejr1OkJ2+CdkRWUICappegbRwOQAWHd43R+4TJr/lG
lKp9ykrsuN4a1sRbo25HhLntS3QV6MGpR1UwBC1fXuHqPeP8lQuMDVtQs2svOhFm
cCdWd/itHD1IliPT7I2dM8GyEq2OJlsugU8VXh6usQVeBZV/NbdqH9+m6gk0Szid
kSP6t9WhMYtP6AMIpX/6xT1ZsyQQSLQOFgi5bdQmSp0xun2OAbq1qBkjoM0qOCnY
k0lVR4x3hNOu2aGLxefF8zdgpZxRMEai8RbJVJW0xk8mCYp6wRYB/o5TYqAAttJV
ai+SEw8kN8RmObnqdCNxW8JEN9Qe22AmMnPJB7GNbxzhV+MlzoaOfuyt2xRZFW8X
X6hxH9RgVyLAdq1RaTBiCVIKxcOLMYR0V/EGmQ9BVLIqAaixDW4BSVJG1Yg+j690
MBteKPnyd4tJYnuu8Mf4Nz2ROVBM9V3T2blhwgUg4loZkDLgaxzky60eyvkFsR16
7IYsTgjw24Vx7EGZ48gKW9ukkPINtWABeplbS+nuI06QNew1L/FhE+jOAofli7+5
S+b82F3GAERNrWa2aGtcqd0YiPBme9Od4wKnPW4bx0V6rt5ad1pGF7d/pN0WtYLu
co5ImTiOlAw56uW+5JFamiyAyZu8BgNf3eR30/y4wD0fh3oPsAxp2HFIci0wWYAz
vyWgl0abUwwgatHqBRL8pCL7X4b+uFtOCZvSeB/3K2fwMO4qEvILz0mBbPxtrv+o
ZLX3HLK6V/yNi/ymkZr59ziPDqi6A+O+cilH+18LHwjH+mvYDl4q8ysek0seS5i9
x2gOYR+k1YNMahl08PeuCxC/bM4W9I7kBZT+OlQu+seVwL/wyex7Wul+4SBdOmQF
r6FbFhbrnsbWJM8ciiyBHPJhrbFgFdVKCoEEo7ssPpILSFRwdiQ8Pci3+jPnyGo+
zVj1WgnvqqD3JGW0C6Vc5YCd6lBgl84AcUTue78lTCdRcrW4/dD0XaEm5WchkxCP
R8ax6n+U3sbZAcwj0N6tsebDuWo9gt6ARAlf235Tx09RvCQKTEjhcV/cvFUh0yOW
H3AV5Bab5GkkIqwUiciPG8FJ/EPvQMaB8gBa0hqQAO58c6Y2PY4j1nfvu/A1liue
xLoP/bL1KL8BAq+j/E3nY2i7x3nsdyL3Jx7Fs3EkAAfskU/SMCpDLZD20x0X+Gl2
ta1VHHmnj5jgVlQPqeTRzmJuFT4ykSry+bSW6J4Z/rwh97wIlmo9oXas8Td/z5RZ
XdEt3uqy4YCMcuz+/FkZHy78R/RcFJaNCE46AjuDLia6a4Ys787LNb8YW43HTF6c
ZFNb9Ji2mQDy+/29bp/gMIdH8gnqgKV45DmTFHIlfDa5JecMRJZ7pHd58+N4dXl+
KY7NCJ5dxfoprQscmeLXfs53UKommUm3P01c/7Msie9qfmEMOkP0WCegqaGZO3dI
ymdGe9Di0QytXC9Q1lRv9WCfWpHgO6eUyhaEJkr6JK90zEef4SQfbyxwvYUnYZn2
aFxbuCUptHdrELEjxTmGiBSGSGk2Vv0bYw6ymjijt7BcU3hlHZ4AOZZRjsaHQYHa
z4cmSiQT9uncRPI0MXnVKMHZ0NX6KcWN14Q/UGeRSOUO+yOmn1k+6iD715TB5FrQ
VhaRYWtVN4dbGKLj+AfWDE8McCCqAA0KobtHDyr7NxnVPSfe+cyHN495zDVRtyTv
R7RKHCqXVsy+NH+gqtHlLAbS+Er7Yi/vW4vdJ2APpKRU4qwXzByifYbuJnAj0t8I
d5hkBocLLxMWGD/JjGr5SCkn3wGSVqui2bkRptdo92SpdKzLXS4cRcUeO/+JvCLb
LNqILl5otnWL6grA6SQKcKoGibOC6eF3XzfaHvnDbG8kbCy5r8EXXi6NRSXNMAxa
w9+UZ0EG2y3CHWHGMRgZxFwc3/vt+4NSEmp/9Dc5YJYP90gWZ7VOMyHVm3pMN5gH
yMtlJ7Vdy+is3w35qU7ypPbYBKb91HFGkGdeH0Z6VavnEpdnmY7EUelVbKkTVxQL
ExQoc4Ucyg54USUjceOOhP2Vc+bAWtrTJsaUKRmzt01jC+b8F2CeV5T6X89zc9Qe
Pa4LyXT5Yed30bfmFFhmkWov/ER5o1MrmNOE4ezw3M4MfctUihypoWVOraRBc7x6
ikmQbYGxm386CVm6WedLh49fukbUYea112YFX1xCtH4ZBbK5PpV3YJSAV0G4/7z/
j/aBA/6EOxdt1E2AnTN3BWS++Apcgdvsglgkm/NNzlJAM4hTT/qxOINhx7OZ0FmS
miHYGcrfmcTBMnXJCrx5RnyII5f6hsd9WoDmCMq3SNMiTaMw9/WhIrNIvO6Uw2Kl
hgYjNGVC7XoJXghtkJwblkcpnVk2hXTQW0rR1Xr/qPE=
`pragma protect end_protected 